/* Machine-generated using Migen */
module top(
	input serial_cts,
	input serial_rts,
	output reg serial_tx,
	input serial_rx,
	input clk200_p,
	input clk200_n,
	input cpu_reset,
	output [15:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output ddram_cs_n,
	output [7:0] ddram_dm,
	inout [63:0] ddram_dq,
	output [7:0] ddram_dqs_p,
	output [7:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash_cs_n,
	inout [3:0] spiflash_dq,
	input eth_clocks_tx,
	output eth_clocks_gtx,
	input eth_clocks_rx,
	output eth_rst_n,
	input eth_int_n,
	input eth_mdio,
	input eth_mdc,
	input eth_rx_dv,
	input eth_rx_er,
	input [7:0] eth_rx_data,
	output reg eth_tx_en,
	output eth_tx_er,
	output reg [7:0] eth_tx_data,
	input eth_col,
	input eth_crs,
	output user_led,
	output user_led_1,
	inout i2c_scl,
	inout i2c_sda,
	output ttl,
	output ttl_1,
	output ttl_2,
	inout ttl_3,
	output ttl_4,
	output ttl_5,
	output ttl_6,
	inout ttl_7,
	output ttl_8,
	output ttl_9,
	output ttl_10,
	inout ttl_11,
	output ttl_12,
	output ttl_13,
	output ttl_14,
	inout ttl_15,
	inout pmt,
	inout pmt_1,
	inout user_sma_gpio_n_33,
	output user_led_2,
	output ams101_dac_ldac,
	inout ams101_dac_clk,
	inout ams101_dac_mosi,
	inout ams101_dac_cs_n,
	output reg la32_p,
	inout spi_clk,
	inout spi_cs_n,
	inout spi_mosi,
	inout spi_miso,
	inout spi_clk_1,
	inout spi_cs_n_1,
	inout spi_mosi_1,
	inout spi_miso_1,
	inout spi_clk_2,
	inout spi_cs_n_2,
	inout spi_mosi_2,
	inout spi_miso_2,
	inout sdcard_spi_33_miso,
	inout sdcard_spi_33_clk,
	inout sdcard_spi_33_mosi,
	inout sdcard_spi_33_cs_n,
	output reg [6:0] dds_a,
	inout [15:0] dds_d,
	output [10:0] dds_sel_n,
	output reg dds_fud,
	output reg dds_wr_n,
	output reg dds_rd_n,
	output dds_rst,
	output reg user_sma_gpio_p_33,
	input user_sma_clock_p,
	input user_sma_clock_n
);

wire [29:0] main_nist_clock_nist_clock_ibus_adr;
wire [31:0] main_nist_clock_nist_clock_ibus_dat_w;
wire [31:0] main_nist_clock_nist_clock_ibus_dat_r;
wire [3:0] main_nist_clock_nist_clock_ibus_sel;
wire main_nist_clock_nist_clock_ibus_cyc;
wire main_nist_clock_nist_clock_ibus_stb;
wire main_nist_clock_nist_clock_ibus_ack;
wire main_nist_clock_nist_clock_ibus_we;
wire [2:0] main_nist_clock_nist_clock_ibus_cti;
wire [1:0] main_nist_clock_nist_clock_ibus_bte;
wire main_nist_clock_nist_clock_ibus_err;
wire [29:0] main_nist_clock_nist_clock_dbus_adr;
wire [31:0] main_nist_clock_nist_clock_dbus_dat_w;
wire [31:0] main_nist_clock_nist_clock_dbus_dat_r;
wire [3:0] main_nist_clock_nist_clock_dbus_sel;
wire main_nist_clock_nist_clock_dbus_cyc;
wire main_nist_clock_nist_clock_dbus_stb;
reg main_nist_clock_nist_clock_dbus_ack;
wire main_nist_clock_nist_clock_dbus_we;
wire [2:0] main_nist_clock_nist_clock_dbus_cti;
wire [1:0] main_nist_clock_nist_clock_dbus_bte;
reg main_nist_clock_nist_clock_dbus_err;
reg [31:0] main_nist_clock_nist_clock_interrupt;
wire [31:0] main_nist_clock_nist_clock_i_adr_o;
wire [31:0] main_nist_clock_nist_clock_d_adr_o;
wire [29:0] main_nist_clock_nist_clock_tmpu_adr;
wire [31:0] main_nist_clock_nist_clock_tmpu_dat_w;
wire [31:0] main_nist_clock_nist_clock_tmpu_dat_r;
wire [3:0] main_nist_clock_nist_clock_tmpu_sel;
wire main_nist_clock_nist_clock_tmpu_cyc;
wire main_nist_clock_nist_clock_tmpu_stb;
wire main_nist_clock_nist_clock_tmpu_ack;
wire main_nist_clock_nist_clock_tmpu_we;
wire [2:0] main_nist_clock_nist_clock_tmpu_cti;
wire [1:0] main_nist_clock_nist_clock_tmpu_bte;
wire main_nist_clock_nist_clock_tmpu_err;
reg main_nist_clock_nist_clock_tmpu_enable_null_storage_full = 1'd0;
wire main_nist_clock_nist_clock_tmpu_enable_null_storage;
reg main_nist_clock_nist_clock_tmpu_enable_null_re = 1'd0;
reg main_nist_clock_nist_clock_tmpu_enable_prog_storage_full = 1'd0;
wire main_nist_clock_nist_clock_tmpu_enable_prog_storage;
reg main_nist_clock_nist_clock_tmpu_enable_prog_re = 1'd0;
reg [29:0] main_nist_clock_nist_clock_tmpu_prog_address_storage_full = 30'd0;
wire [17:0] main_nist_clock_nist_clock_tmpu_prog_address_storage;
reg main_nist_clock_nist_clock_tmpu_prog_address_re = 1'd0;
reg main_nist_clock_nist_clock_tmpu_error = 1'd0;
wire [29:0] main_nist_clock_nist_clock_sram_bus_adr;
wire [31:0] main_nist_clock_nist_clock_sram_bus_dat_w;
wire [31:0] main_nist_clock_nist_clock_sram_bus_dat_r;
wire [3:0] main_nist_clock_nist_clock_sram_bus_sel;
wire main_nist_clock_nist_clock_sram_bus_cyc;
wire main_nist_clock_nist_clock_sram_bus_stb;
reg main_nist_clock_nist_clock_sram_bus_ack = 1'd0;
wire main_nist_clock_nist_clock_sram_bus_we;
wire [2:0] main_nist_clock_nist_clock_sram_bus_cti;
wire [1:0] main_nist_clock_nist_clock_sram_bus_bte;
reg main_nist_clock_nist_clock_sram_bus_err = 1'd0;
wire [10:0] main_nist_clock_nist_clock_sram_adr;
wire [31:0] main_nist_clock_nist_clock_sram_dat_r;
reg [3:0] main_nist_clock_nist_clock_sram_we;
wire [31:0] main_nist_clock_nist_clock_sram_dat_w;
reg [13:0] main_nist_clock_nist_clock_interface_adr = 14'd0;
reg main_nist_clock_nist_clock_interface_we = 1'd0;
reg [7:0] main_nist_clock_nist_clock_interface_dat_w = 8'd0;
wire [7:0] main_nist_clock_nist_clock_interface_dat_r;
wire [29:0] main_nist_clock_nist_clock_bus_wishbone_adr;
wire [31:0] main_nist_clock_nist_clock_bus_wishbone_dat_w;
reg [31:0] main_nist_clock_nist_clock_bus_wishbone_dat_r = 32'd0;
wire [3:0] main_nist_clock_nist_clock_bus_wishbone_sel;
wire main_nist_clock_nist_clock_bus_wishbone_cyc;
wire main_nist_clock_nist_clock_bus_wishbone_stb;
reg main_nist_clock_nist_clock_bus_wishbone_ack = 1'd0;
wire main_nist_clock_nist_clock_bus_wishbone_we;
wire [2:0] main_nist_clock_nist_clock_bus_wishbone_cti;
wire [1:0] main_nist_clock_nist_clock_bus_wishbone_bte;
reg main_nist_clock_nist_clock_bus_wishbone_err = 1'd0;
reg [1:0] main_nist_clock_nist_clock_counter = 2'd0;
reg [31:0] main_nist_clock_nist_clock_uart_phy_storage_full = 32'd3958241;
wire [31:0] main_nist_clock_nist_clock_uart_phy_storage;
reg main_nist_clock_nist_clock_uart_phy_re = 1'd0;
wire main_nist_clock_nist_clock_uart_phy_sink_stb;
reg main_nist_clock_nist_clock_uart_phy_sink_ack = 1'd0;
wire main_nist_clock_nist_clock_uart_phy_sink_eop;
wire [7:0] main_nist_clock_nist_clock_uart_phy_sink_payload_data;
reg main_nist_clock_nist_clock_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] main_nist_clock_nist_clock_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] main_nist_clock_nist_clock_uart_phy_tx_reg = 8'd0;
reg [3:0] main_nist_clock_nist_clock_uart_phy_tx_bitcount = 4'd0;
reg main_nist_clock_nist_clock_uart_phy_tx_busy = 1'd0;
reg main_nist_clock_nist_clock_uart_phy_source_stb = 1'd0;
wire main_nist_clock_nist_clock_uart_phy_source_ack;
reg main_nist_clock_nist_clock_uart_phy_source_eop = 1'd0;
reg [7:0] main_nist_clock_nist_clock_uart_phy_source_payload_data = 8'd0;
reg main_nist_clock_nist_clock_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] main_nist_clock_nist_clock_uart_phy_phase_accumulator_rx = 32'd0;
wire main_nist_clock_nist_clock_uart_phy_rx;
reg main_nist_clock_nist_clock_uart_phy_rx_r = 1'd0;
reg [7:0] main_nist_clock_nist_clock_uart_phy_rx_reg = 8'd0;
reg [3:0] main_nist_clock_nist_clock_uart_phy_rx_bitcount = 4'd0;
reg main_nist_clock_nist_clock_uart_phy_rx_busy = 1'd0;
wire main_nist_clock_nist_clock_uart_rxtx_re;
wire [7:0] main_nist_clock_nist_clock_uart_rxtx_r;
wire [7:0] main_nist_clock_nist_clock_uart_rxtx_w;
wire main_nist_clock_nist_clock_uart_txfull_status;
wire main_nist_clock_nist_clock_uart_rxempty_status;
wire main_nist_clock_nist_clock_uart_irq;
wire main_nist_clock_nist_clock_uart_tx_status;
reg main_nist_clock_nist_clock_uart_tx_pending = 1'd0;
wire main_nist_clock_nist_clock_uart_tx_trigger;
reg main_nist_clock_nist_clock_uart_tx_clear;
reg main_nist_clock_nist_clock_uart_tx_old_trigger = 1'd0;
wire main_nist_clock_nist_clock_uart_rx_status;
reg main_nist_clock_nist_clock_uart_rx_pending = 1'd0;
wire main_nist_clock_nist_clock_uart_rx_trigger;
reg main_nist_clock_nist_clock_uart_rx_clear;
reg main_nist_clock_nist_clock_uart_rx_old_trigger = 1'd0;
wire main_nist_clock_nist_clock_uart_status_re;
wire [1:0] main_nist_clock_nist_clock_uart_status_r;
reg [1:0] main_nist_clock_nist_clock_uart_status_w;
wire main_nist_clock_nist_clock_uart_pending_re;
wire [1:0] main_nist_clock_nist_clock_uart_pending_r;
reg [1:0] main_nist_clock_nist_clock_uart_pending_w;
reg [1:0] main_nist_clock_nist_clock_uart_storage_full = 2'd0;
wire [1:0] main_nist_clock_nist_clock_uart_storage;
reg main_nist_clock_nist_clock_uart_re = 1'd0;
wire main_nist_clock_nist_clock_uart_tx_fifo_sink_stb;
wire main_nist_clock_nist_clock_uart_tx_fifo_sink_ack;
reg main_nist_clock_nist_clock_uart_tx_fifo_sink_eop = 1'd0;
wire [7:0] main_nist_clock_nist_clock_uart_tx_fifo_sink_payload_data;
wire main_nist_clock_nist_clock_uart_tx_fifo_source_stb;
wire main_nist_clock_nist_clock_uart_tx_fifo_source_ack;
wire main_nist_clock_nist_clock_uart_tx_fifo_source_eop;
wire [7:0] main_nist_clock_nist_clock_uart_tx_fifo_source_payload_data;
wire main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_we;
wire main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable;
wire main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_re;
wire main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_readable;
wire [8:0] main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_din;
wire [8:0] main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_dout;
reg [4:0] main_nist_clock_nist_clock_uart_tx_fifo_level = 5'd0;
reg main_nist_clock_nist_clock_uart_tx_fifo_replace = 1'd0;
reg [3:0] main_nist_clock_nist_clock_uart_tx_fifo_produce = 4'd0;
reg [3:0] main_nist_clock_nist_clock_uart_tx_fifo_consume = 4'd0;
reg [3:0] main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr;
wire [8:0] main_nist_clock_nist_clock_uart_tx_fifo_wrport_dat_r;
wire main_nist_clock_nist_clock_uart_tx_fifo_wrport_we;
wire [8:0] main_nist_clock_nist_clock_uart_tx_fifo_wrport_dat_w;
wire main_nist_clock_nist_clock_uart_tx_fifo_do_read;
wire [3:0] main_nist_clock_nist_clock_uart_tx_fifo_rdport_adr;
wire [8:0] main_nist_clock_nist_clock_uart_tx_fifo_rdport_dat_r;
wire [7:0] main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_payload_data;
wire main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_eop;
wire [7:0] main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_payload_data;
wire main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_eop;
wire main_nist_clock_nist_clock_uart_rx_fifo_sink_stb;
wire main_nist_clock_nist_clock_uart_rx_fifo_sink_ack;
wire main_nist_clock_nist_clock_uart_rx_fifo_sink_eop;
wire [7:0] main_nist_clock_nist_clock_uart_rx_fifo_sink_payload_data;
wire main_nist_clock_nist_clock_uart_rx_fifo_source_stb;
wire main_nist_clock_nist_clock_uart_rx_fifo_source_ack;
wire main_nist_clock_nist_clock_uart_rx_fifo_source_eop;
wire [7:0] main_nist_clock_nist_clock_uart_rx_fifo_source_payload_data;
wire main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_we;
wire main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable;
wire main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_re;
wire main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_readable;
wire [8:0] main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_din;
wire [8:0] main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_dout;
reg [4:0] main_nist_clock_nist_clock_uart_rx_fifo_level = 5'd0;
reg main_nist_clock_nist_clock_uart_rx_fifo_replace = 1'd0;
reg [3:0] main_nist_clock_nist_clock_uart_rx_fifo_produce = 4'd0;
reg [3:0] main_nist_clock_nist_clock_uart_rx_fifo_consume = 4'd0;
reg [3:0] main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr;
wire [8:0] main_nist_clock_nist_clock_uart_rx_fifo_wrport_dat_r;
wire main_nist_clock_nist_clock_uart_rx_fifo_wrport_we;
wire [8:0] main_nist_clock_nist_clock_uart_rx_fifo_wrport_dat_w;
wire main_nist_clock_nist_clock_uart_rx_fifo_do_read;
wire [3:0] main_nist_clock_nist_clock_uart_rx_fifo_rdport_adr;
wire [8:0] main_nist_clock_nist_clock_uart_rx_fifo_rdport_dat_r;
wire [7:0] main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_payload_data;
wire main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_eop;
wire [7:0] main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_payload_data;
wire main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_eop;
reg [63:0] main_nist_clock_nist_clock_timer0_load_storage_full = 64'd0;
wire [63:0] main_nist_clock_nist_clock_timer0_load_storage;
reg main_nist_clock_nist_clock_timer0_load_re = 1'd0;
reg [63:0] main_nist_clock_nist_clock_timer0_reload_storage_full = 64'd0;
wire [63:0] main_nist_clock_nist_clock_timer0_reload_storage;
reg main_nist_clock_nist_clock_timer0_reload_re = 1'd0;
reg main_nist_clock_nist_clock_timer0_en_storage_full = 1'd0;
wire main_nist_clock_nist_clock_timer0_en_storage;
reg main_nist_clock_nist_clock_timer0_en_re = 1'd0;
wire main_nist_clock_nist_clock_timer0_update_value_re;
wire main_nist_clock_nist_clock_timer0_update_value_r;
reg main_nist_clock_nist_clock_timer0_update_value_w = 1'd0;
reg [63:0] main_nist_clock_nist_clock_timer0_value_status = 64'd0;
wire main_nist_clock_nist_clock_timer0_irq;
wire main_nist_clock_nist_clock_timer0_zero_status;
reg main_nist_clock_nist_clock_timer0_zero_pending = 1'd0;
wire main_nist_clock_nist_clock_timer0_zero_trigger;
reg main_nist_clock_nist_clock_timer0_zero_clear;
reg main_nist_clock_nist_clock_timer0_zero_old_trigger = 1'd0;
wire main_nist_clock_nist_clock_timer0_eventmanager_status_re;
wire main_nist_clock_nist_clock_timer0_eventmanager_status_r;
wire main_nist_clock_nist_clock_timer0_eventmanager_status_w;
wire main_nist_clock_nist_clock_timer0_eventmanager_pending_re;
wire main_nist_clock_nist_clock_timer0_eventmanager_pending_r;
wire main_nist_clock_nist_clock_timer0_eventmanager_pending_w;
reg main_nist_clock_nist_clock_timer0_eventmanager_storage_full = 1'd0;
wire main_nist_clock_nist_clock_timer0_eventmanager_storage;
reg main_nist_clock_nist_clock_timer0_eventmanager_re = 1'd0;
reg [63:0] main_nist_clock_nist_clock_timer0_value = 64'd0;
wire [29:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr;
wire [31:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_w;
reg [31:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r;
wire [3:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel;
wire main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cyc;
wire main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_stb;
reg main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack;
wire main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_we;
wire [2:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cti;
wire [1:0] main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_bte;
reg main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire clk200_clk;
wire clk200_rst;
wire main_nist_clock_clk200_se;
wire main_nist_clock_pll_locked;
wire main_nist_clock_pll_fb;
wire main_nist_clock_pll_sys;
wire main_nist_clock_pll_sys4x;
wire main_nist_clock_pll_clk200;
reg [3:0] main_nist_clock_reset_counter = 4'd15;
reg main_nist_clock_ic_reset = 1'd1;
reg main_nist_clock_ddrphy_wlevel_en_storage_full = 1'd0;
wire main_nist_clock_ddrphy_wlevel_en_storage;
reg main_nist_clock_ddrphy_wlevel_en_re = 1'd0;
wire main_nist_clock_ddrphy_wlevel_strobe_re;
wire main_nist_clock_ddrphy_wlevel_strobe_r;
reg main_nist_clock_ddrphy_wlevel_strobe_w = 1'd0;
reg [7:0] main_nist_clock_ddrphy_dly_sel_storage_full = 8'd0;
wire [7:0] main_nist_clock_ddrphy_dly_sel_storage;
reg main_nist_clock_ddrphy_dly_sel_re = 1'd0;
wire main_nist_clock_ddrphy_rdly_dq_rst_re;
wire main_nist_clock_ddrphy_rdly_dq_rst_r;
reg main_nist_clock_ddrphy_rdly_dq_rst_w = 1'd0;
wire main_nist_clock_ddrphy_rdly_dq_inc_re;
wire main_nist_clock_ddrphy_rdly_dq_inc_r;
reg main_nist_clock_ddrphy_rdly_dq_inc_w = 1'd0;
wire main_nist_clock_ddrphy_rdly_dq_bitslip_re;
wire main_nist_clock_ddrphy_rdly_dq_bitslip_r;
reg main_nist_clock_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire main_nist_clock_ddrphy_wdly_dq_rst_re;
wire main_nist_clock_ddrphy_wdly_dq_rst_r;
reg main_nist_clock_ddrphy_wdly_dq_rst_w = 1'd0;
wire main_nist_clock_ddrphy_wdly_dq_inc_re;
wire main_nist_clock_ddrphy_wdly_dq_inc_r;
reg main_nist_clock_ddrphy_wdly_dq_inc_w = 1'd0;
wire main_nist_clock_ddrphy_wdly_dqs_rst_re;
wire main_nist_clock_ddrphy_wdly_dqs_rst_r;
reg main_nist_clock_ddrphy_wdly_dqs_rst_w = 1'd0;
wire main_nist_clock_ddrphy_wdly_dqs_inc_re;
wire main_nist_clock_ddrphy_wdly_dqs_inc_r;
reg main_nist_clock_ddrphy_wdly_dqs_inc_w = 1'd0;
wire [15:0] main_nist_clock_ddrphy_dfi_p0_address;
wire [2:0] main_nist_clock_ddrphy_dfi_p0_bank;
wire main_nist_clock_ddrphy_dfi_p0_cas_n;
wire main_nist_clock_ddrphy_dfi_p0_cs_n;
wire main_nist_clock_ddrphy_dfi_p0_ras_n;
wire main_nist_clock_ddrphy_dfi_p0_we_n;
wire main_nist_clock_ddrphy_dfi_p0_cke;
wire main_nist_clock_ddrphy_dfi_p0_odt;
wire main_nist_clock_ddrphy_dfi_p0_reset_n;
wire [127:0] main_nist_clock_ddrphy_dfi_p0_wrdata;
wire main_nist_clock_ddrphy_dfi_p0_wrdata_en;
wire [15:0] main_nist_clock_ddrphy_dfi_p0_wrdata_mask;
wire main_nist_clock_ddrphy_dfi_p0_rddata_en;
wire [127:0] main_nist_clock_ddrphy_dfi_p0_rddata;
reg main_nist_clock_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [15:0] main_nist_clock_ddrphy_dfi_p1_address;
wire [2:0] main_nist_clock_ddrphy_dfi_p1_bank;
wire main_nist_clock_ddrphy_dfi_p1_cas_n;
wire main_nist_clock_ddrphy_dfi_p1_cs_n;
wire main_nist_clock_ddrphy_dfi_p1_ras_n;
wire main_nist_clock_ddrphy_dfi_p1_we_n;
wire main_nist_clock_ddrphy_dfi_p1_cke;
wire main_nist_clock_ddrphy_dfi_p1_odt;
wire main_nist_clock_ddrphy_dfi_p1_reset_n;
wire [127:0] main_nist_clock_ddrphy_dfi_p1_wrdata;
wire main_nist_clock_ddrphy_dfi_p1_wrdata_en;
wire [15:0] main_nist_clock_ddrphy_dfi_p1_wrdata_mask;
wire main_nist_clock_ddrphy_dfi_p1_rddata_en;
wire [127:0] main_nist_clock_ddrphy_dfi_p1_rddata;
reg main_nist_clock_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [15:0] main_nist_clock_ddrphy_dfi_p2_address;
wire [2:0] main_nist_clock_ddrphy_dfi_p2_bank;
wire main_nist_clock_ddrphy_dfi_p2_cas_n;
wire main_nist_clock_ddrphy_dfi_p2_cs_n;
wire main_nist_clock_ddrphy_dfi_p2_ras_n;
wire main_nist_clock_ddrphy_dfi_p2_we_n;
wire main_nist_clock_ddrphy_dfi_p2_cke;
wire main_nist_clock_ddrphy_dfi_p2_odt;
wire main_nist_clock_ddrphy_dfi_p2_reset_n;
wire [127:0] main_nist_clock_ddrphy_dfi_p2_wrdata;
wire main_nist_clock_ddrphy_dfi_p2_wrdata_en;
wire [15:0] main_nist_clock_ddrphy_dfi_p2_wrdata_mask;
wire main_nist_clock_ddrphy_dfi_p2_rddata_en;
wire [127:0] main_nist_clock_ddrphy_dfi_p2_rddata;
reg main_nist_clock_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [15:0] main_nist_clock_ddrphy_dfi_p3_address;
wire [2:0] main_nist_clock_ddrphy_dfi_p3_bank;
wire main_nist_clock_ddrphy_dfi_p3_cas_n;
wire main_nist_clock_ddrphy_dfi_p3_cs_n;
wire main_nist_clock_ddrphy_dfi_p3_ras_n;
wire main_nist_clock_ddrphy_dfi_p3_we_n;
wire main_nist_clock_ddrphy_dfi_p3_cke;
wire main_nist_clock_ddrphy_dfi_p3_odt;
wire main_nist_clock_ddrphy_dfi_p3_reset_n;
wire [127:0] main_nist_clock_ddrphy_dfi_p3_wrdata;
wire main_nist_clock_ddrphy_dfi_p3_wrdata_en;
wire [15:0] main_nist_clock_ddrphy_dfi_p3_wrdata_mask;
wire main_nist_clock_ddrphy_dfi_p3_rddata_en;
wire [127:0] main_nist_clock_ddrphy_dfi_p3_rddata;
reg main_nist_clock_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire main_nist_clock_ddrphy_sd_clk_se;
reg main_nist_clock_ddrphy_oe_dqs = 1'd0;
reg [7:0] main_nist_clock_ddrphy_dqs_serdes_pattern;
wire main_nist_clock_ddrphy_dm_o_nodelay0;
wire main_nist_clock_ddrphy_dqs_nodelay0;
wire main_nist_clock_ddrphy_dqs_delayed0;
wire main_nist_clock_ddrphy_dqs_t0;
wire main_nist_clock_ddrphy_dm_o_nodelay1;
wire main_nist_clock_ddrphy_dqs_nodelay1;
wire main_nist_clock_ddrphy_dqs_delayed1;
wire main_nist_clock_ddrphy_dqs_t1;
wire main_nist_clock_ddrphy_dm_o_nodelay2;
wire main_nist_clock_ddrphy_dqs_nodelay2;
wire main_nist_clock_ddrphy_dqs_delayed2;
wire main_nist_clock_ddrphy_dqs_t2;
wire main_nist_clock_ddrphy_dm_o_nodelay3;
wire main_nist_clock_ddrphy_dqs_nodelay3;
wire main_nist_clock_ddrphy_dqs_delayed3;
wire main_nist_clock_ddrphy_dqs_t3;
wire main_nist_clock_ddrphy_dm_o_nodelay4;
wire main_nist_clock_ddrphy_dqs_nodelay4;
wire main_nist_clock_ddrphy_dqs_delayed4;
wire main_nist_clock_ddrphy_dqs_t4;
wire main_nist_clock_ddrphy_dm_o_nodelay5;
wire main_nist_clock_ddrphy_dqs_nodelay5;
wire main_nist_clock_ddrphy_dqs_delayed5;
wire main_nist_clock_ddrphy_dqs_t5;
wire main_nist_clock_ddrphy_dm_o_nodelay6;
wire main_nist_clock_ddrphy_dqs_nodelay6;
wire main_nist_clock_ddrphy_dqs_delayed6;
wire main_nist_clock_ddrphy_dqs_t6;
wire main_nist_clock_ddrphy_dm_o_nodelay7;
wire main_nist_clock_ddrphy_dqs_nodelay7;
wire main_nist_clock_ddrphy_dqs_delayed7;
wire main_nist_clock_ddrphy_dqs_t7;
reg main_nist_clock_ddrphy_oe_dq = 1'd0;
wire main_nist_clock_ddrphy_dq_o_nodelay0;
wire main_nist_clock_ddrphy_dq_o_delayed0;
wire main_nist_clock_ddrphy_dq_i_nodelay0;
wire main_nist_clock_ddrphy_dq_i_delayed0;
wire main_nist_clock_ddrphy_dq_t0;
wire main_nist_clock_ddrphy_dq_o_nodelay1;
wire main_nist_clock_ddrphy_dq_o_delayed1;
wire main_nist_clock_ddrphy_dq_i_nodelay1;
wire main_nist_clock_ddrphy_dq_i_delayed1;
wire main_nist_clock_ddrphy_dq_t1;
wire main_nist_clock_ddrphy_dq_o_nodelay2;
wire main_nist_clock_ddrphy_dq_o_delayed2;
wire main_nist_clock_ddrphy_dq_i_nodelay2;
wire main_nist_clock_ddrphy_dq_i_delayed2;
wire main_nist_clock_ddrphy_dq_t2;
wire main_nist_clock_ddrphy_dq_o_nodelay3;
wire main_nist_clock_ddrphy_dq_o_delayed3;
wire main_nist_clock_ddrphy_dq_i_nodelay3;
wire main_nist_clock_ddrphy_dq_i_delayed3;
wire main_nist_clock_ddrphy_dq_t3;
wire main_nist_clock_ddrphy_dq_o_nodelay4;
wire main_nist_clock_ddrphy_dq_o_delayed4;
wire main_nist_clock_ddrphy_dq_i_nodelay4;
wire main_nist_clock_ddrphy_dq_i_delayed4;
wire main_nist_clock_ddrphy_dq_t4;
wire main_nist_clock_ddrphy_dq_o_nodelay5;
wire main_nist_clock_ddrphy_dq_o_delayed5;
wire main_nist_clock_ddrphy_dq_i_nodelay5;
wire main_nist_clock_ddrphy_dq_i_delayed5;
wire main_nist_clock_ddrphy_dq_t5;
wire main_nist_clock_ddrphy_dq_o_nodelay6;
wire main_nist_clock_ddrphy_dq_o_delayed6;
wire main_nist_clock_ddrphy_dq_i_nodelay6;
wire main_nist_clock_ddrphy_dq_i_delayed6;
wire main_nist_clock_ddrphy_dq_t6;
wire main_nist_clock_ddrphy_dq_o_nodelay7;
wire main_nist_clock_ddrphy_dq_o_delayed7;
wire main_nist_clock_ddrphy_dq_i_nodelay7;
wire main_nist_clock_ddrphy_dq_i_delayed7;
wire main_nist_clock_ddrphy_dq_t7;
wire main_nist_clock_ddrphy_dq_o_nodelay8;
wire main_nist_clock_ddrphy_dq_o_delayed8;
wire main_nist_clock_ddrphy_dq_i_nodelay8;
wire main_nist_clock_ddrphy_dq_i_delayed8;
wire main_nist_clock_ddrphy_dq_t8;
wire main_nist_clock_ddrphy_dq_o_nodelay9;
wire main_nist_clock_ddrphy_dq_o_delayed9;
wire main_nist_clock_ddrphy_dq_i_nodelay9;
wire main_nist_clock_ddrphy_dq_i_delayed9;
wire main_nist_clock_ddrphy_dq_t9;
wire main_nist_clock_ddrphy_dq_o_nodelay10;
wire main_nist_clock_ddrphy_dq_o_delayed10;
wire main_nist_clock_ddrphy_dq_i_nodelay10;
wire main_nist_clock_ddrphy_dq_i_delayed10;
wire main_nist_clock_ddrphy_dq_t10;
wire main_nist_clock_ddrphy_dq_o_nodelay11;
wire main_nist_clock_ddrphy_dq_o_delayed11;
wire main_nist_clock_ddrphy_dq_i_nodelay11;
wire main_nist_clock_ddrphy_dq_i_delayed11;
wire main_nist_clock_ddrphy_dq_t11;
wire main_nist_clock_ddrphy_dq_o_nodelay12;
wire main_nist_clock_ddrphy_dq_o_delayed12;
wire main_nist_clock_ddrphy_dq_i_nodelay12;
wire main_nist_clock_ddrphy_dq_i_delayed12;
wire main_nist_clock_ddrphy_dq_t12;
wire main_nist_clock_ddrphy_dq_o_nodelay13;
wire main_nist_clock_ddrphy_dq_o_delayed13;
wire main_nist_clock_ddrphy_dq_i_nodelay13;
wire main_nist_clock_ddrphy_dq_i_delayed13;
wire main_nist_clock_ddrphy_dq_t13;
wire main_nist_clock_ddrphy_dq_o_nodelay14;
wire main_nist_clock_ddrphy_dq_o_delayed14;
wire main_nist_clock_ddrphy_dq_i_nodelay14;
wire main_nist_clock_ddrphy_dq_i_delayed14;
wire main_nist_clock_ddrphy_dq_t14;
wire main_nist_clock_ddrphy_dq_o_nodelay15;
wire main_nist_clock_ddrphy_dq_o_delayed15;
wire main_nist_clock_ddrphy_dq_i_nodelay15;
wire main_nist_clock_ddrphy_dq_i_delayed15;
wire main_nist_clock_ddrphy_dq_t15;
wire main_nist_clock_ddrphy_dq_o_nodelay16;
wire main_nist_clock_ddrphy_dq_o_delayed16;
wire main_nist_clock_ddrphy_dq_i_nodelay16;
wire main_nist_clock_ddrphy_dq_i_delayed16;
wire main_nist_clock_ddrphy_dq_t16;
wire main_nist_clock_ddrphy_dq_o_nodelay17;
wire main_nist_clock_ddrphy_dq_o_delayed17;
wire main_nist_clock_ddrphy_dq_i_nodelay17;
wire main_nist_clock_ddrphy_dq_i_delayed17;
wire main_nist_clock_ddrphy_dq_t17;
wire main_nist_clock_ddrphy_dq_o_nodelay18;
wire main_nist_clock_ddrphy_dq_o_delayed18;
wire main_nist_clock_ddrphy_dq_i_nodelay18;
wire main_nist_clock_ddrphy_dq_i_delayed18;
wire main_nist_clock_ddrphy_dq_t18;
wire main_nist_clock_ddrphy_dq_o_nodelay19;
wire main_nist_clock_ddrphy_dq_o_delayed19;
wire main_nist_clock_ddrphy_dq_i_nodelay19;
wire main_nist_clock_ddrphy_dq_i_delayed19;
wire main_nist_clock_ddrphy_dq_t19;
wire main_nist_clock_ddrphy_dq_o_nodelay20;
wire main_nist_clock_ddrphy_dq_o_delayed20;
wire main_nist_clock_ddrphy_dq_i_nodelay20;
wire main_nist_clock_ddrphy_dq_i_delayed20;
wire main_nist_clock_ddrphy_dq_t20;
wire main_nist_clock_ddrphy_dq_o_nodelay21;
wire main_nist_clock_ddrphy_dq_o_delayed21;
wire main_nist_clock_ddrphy_dq_i_nodelay21;
wire main_nist_clock_ddrphy_dq_i_delayed21;
wire main_nist_clock_ddrphy_dq_t21;
wire main_nist_clock_ddrphy_dq_o_nodelay22;
wire main_nist_clock_ddrphy_dq_o_delayed22;
wire main_nist_clock_ddrphy_dq_i_nodelay22;
wire main_nist_clock_ddrphy_dq_i_delayed22;
wire main_nist_clock_ddrphy_dq_t22;
wire main_nist_clock_ddrphy_dq_o_nodelay23;
wire main_nist_clock_ddrphy_dq_o_delayed23;
wire main_nist_clock_ddrphy_dq_i_nodelay23;
wire main_nist_clock_ddrphy_dq_i_delayed23;
wire main_nist_clock_ddrphy_dq_t23;
wire main_nist_clock_ddrphy_dq_o_nodelay24;
wire main_nist_clock_ddrphy_dq_o_delayed24;
wire main_nist_clock_ddrphy_dq_i_nodelay24;
wire main_nist_clock_ddrphy_dq_i_delayed24;
wire main_nist_clock_ddrphy_dq_t24;
wire main_nist_clock_ddrphy_dq_o_nodelay25;
wire main_nist_clock_ddrphy_dq_o_delayed25;
wire main_nist_clock_ddrphy_dq_i_nodelay25;
wire main_nist_clock_ddrphy_dq_i_delayed25;
wire main_nist_clock_ddrphy_dq_t25;
wire main_nist_clock_ddrphy_dq_o_nodelay26;
wire main_nist_clock_ddrphy_dq_o_delayed26;
wire main_nist_clock_ddrphy_dq_i_nodelay26;
wire main_nist_clock_ddrphy_dq_i_delayed26;
wire main_nist_clock_ddrphy_dq_t26;
wire main_nist_clock_ddrphy_dq_o_nodelay27;
wire main_nist_clock_ddrphy_dq_o_delayed27;
wire main_nist_clock_ddrphy_dq_i_nodelay27;
wire main_nist_clock_ddrphy_dq_i_delayed27;
wire main_nist_clock_ddrphy_dq_t27;
wire main_nist_clock_ddrphy_dq_o_nodelay28;
wire main_nist_clock_ddrphy_dq_o_delayed28;
wire main_nist_clock_ddrphy_dq_i_nodelay28;
wire main_nist_clock_ddrphy_dq_i_delayed28;
wire main_nist_clock_ddrphy_dq_t28;
wire main_nist_clock_ddrphy_dq_o_nodelay29;
wire main_nist_clock_ddrphy_dq_o_delayed29;
wire main_nist_clock_ddrphy_dq_i_nodelay29;
wire main_nist_clock_ddrphy_dq_i_delayed29;
wire main_nist_clock_ddrphy_dq_t29;
wire main_nist_clock_ddrphy_dq_o_nodelay30;
wire main_nist_clock_ddrphy_dq_o_delayed30;
wire main_nist_clock_ddrphy_dq_i_nodelay30;
wire main_nist_clock_ddrphy_dq_i_delayed30;
wire main_nist_clock_ddrphy_dq_t30;
wire main_nist_clock_ddrphy_dq_o_nodelay31;
wire main_nist_clock_ddrphy_dq_o_delayed31;
wire main_nist_clock_ddrphy_dq_i_nodelay31;
wire main_nist_clock_ddrphy_dq_i_delayed31;
wire main_nist_clock_ddrphy_dq_t31;
wire main_nist_clock_ddrphy_dq_o_nodelay32;
wire main_nist_clock_ddrphy_dq_o_delayed32;
wire main_nist_clock_ddrphy_dq_i_nodelay32;
wire main_nist_clock_ddrphy_dq_i_delayed32;
wire main_nist_clock_ddrphy_dq_t32;
wire main_nist_clock_ddrphy_dq_o_nodelay33;
wire main_nist_clock_ddrphy_dq_o_delayed33;
wire main_nist_clock_ddrphy_dq_i_nodelay33;
wire main_nist_clock_ddrphy_dq_i_delayed33;
wire main_nist_clock_ddrphy_dq_t33;
wire main_nist_clock_ddrphy_dq_o_nodelay34;
wire main_nist_clock_ddrphy_dq_o_delayed34;
wire main_nist_clock_ddrphy_dq_i_nodelay34;
wire main_nist_clock_ddrphy_dq_i_delayed34;
wire main_nist_clock_ddrphy_dq_t34;
wire main_nist_clock_ddrphy_dq_o_nodelay35;
wire main_nist_clock_ddrphy_dq_o_delayed35;
wire main_nist_clock_ddrphy_dq_i_nodelay35;
wire main_nist_clock_ddrphy_dq_i_delayed35;
wire main_nist_clock_ddrphy_dq_t35;
wire main_nist_clock_ddrphy_dq_o_nodelay36;
wire main_nist_clock_ddrphy_dq_o_delayed36;
wire main_nist_clock_ddrphy_dq_i_nodelay36;
wire main_nist_clock_ddrphy_dq_i_delayed36;
wire main_nist_clock_ddrphy_dq_t36;
wire main_nist_clock_ddrphy_dq_o_nodelay37;
wire main_nist_clock_ddrphy_dq_o_delayed37;
wire main_nist_clock_ddrphy_dq_i_nodelay37;
wire main_nist_clock_ddrphy_dq_i_delayed37;
wire main_nist_clock_ddrphy_dq_t37;
wire main_nist_clock_ddrphy_dq_o_nodelay38;
wire main_nist_clock_ddrphy_dq_o_delayed38;
wire main_nist_clock_ddrphy_dq_i_nodelay38;
wire main_nist_clock_ddrphy_dq_i_delayed38;
wire main_nist_clock_ddrphy_dq_t38;
wire main_nist_clock_ddrphy_dq_o_nodelay39;
wire main_nist_clock_ddrphy_dq_o_delayed39;
wire main_nist_clock_ddrphy_dq_i_nodelay39;
wire main_nist_clock_ddrphy_dq_i_delayed39;
wire main_nist_clock_ddrphy_dq_t39;
wire main_nist_clock_ddrphy_dq_o_nodelay40;
wire main_nist_clock_ddrphy_dq_o_delayed40;
wire main_nist_clock_ddrphy_dq_i_nodelay40;
wire main_nist_clock_ddrphy_dq_i_delayed40;
wire main_nist_clock_ddrphy_dq_t40;
wire main_nist_clock_ddrphy_dq_o_nodelay41;
wire main_nist_clock_ddrphy_dq_o_delayed41;
wire main_nist_clock_ddrphy_dq_i_nodelay41;
wire main_nist_clock_ddrphy_dq_i_delayed41;
wire main_nist_clock_ddrphy_dq_t41;
wire main_nist_clock_ddrphy_dq_o_nodelay42;
wire main_nist_clock_ddrphy_dq_o_delayed42;
wire main_nist_clock_ddrphy_dq_i_nodelay42;
wire main_nist_clock_ddrphy_dq_i_delayed42;
wire main_nist_clock_ddrphy_dq_t42;
wire main_nist_clock_ddrphy_dq_o_nodelay43;
wire main_nist_clock_ddrphy_dq_o_delayed43;
wire main_nist_clock_ddrphy_dq_i_nodelay43;
wire main_nist_clock_ddrphy_dq_i_delayed43;
wire main_nist_clock_ddrphy_dq_t43;
wire main_nist_clock_ddrphy_dq_o_nodelay44;
wire main_nist_clock_ddrphy_dq_o_delayed44;
wire main_nist_clock_ddrphy_dq_i_nodelay44;
wire main_nist_clock_ddrphy_dq_i_delayed44;
wire main_nist_clock_ddrphy_dq_t44;
wire main_nist_clock_ddrphy_dq_o_nodelay45;
wire main_nist_clock_ddrphy_dq_o_delayed45;
wire main_nist_clock_ddrphy_dq_i_nodelay45;
wire main_nist_clock_ddrphy_dq_i_delayed45;
wire main_nist_clock_ddrphy_dq_t45;
wire main_nist_clock_ddrphy_dq_o_nodelay46;
wire main_nist_clock_ddrphy_dq_o_delayed46;
wire main_nist_clock_ddrphy_dq_i_nodelay46;
wire main_nist_clock_ddrphy_dq_i_delayed46;
wire main_nist_clock_ddrphy_dq_t46;
wire main_nist_clock_ddrphy_dq_o_nodelay47;
wire main_nist_clock_ddrphy_dq_o_delayed47;
wire main_nist_clock_ddrphy_dq_i_nodelay47;
wire main_nist_clock_ddrphy_dq_i_delayed47;
wire main_nist_clock_ddrphy_dq_t47;
wire main_nist_clock_ddrphy_dq_o_nodelay48;
wire main_nist_clock_ddrphy_dq_o_delayed48;
wire main_nist_clock_ddrphy_dq_i_nodelay48;
wire main_nist_clock_ddrphy_dq_i_delayed48;
wire main_nist_clock_ddrphy_dq_t48;
wire main_nist_clock_ddrphy_dq_o_nodelay49;
wire main_nist_clock_ddrphy_dq_o_delayed49;
wire main_nist_clock_ddrphy_dq_i_nodelay49;
wire main_nist_clock_ddrphy_dq_i_delayed49;
wire main_nist_clock_ddrphy_dq_t49;
wire main_nist_clock_ddrphy_dq_o_nodelay50;
wire main_nist_clock_ddrphy_dq_o_delayed50;
wire main_nist_clock_ddrphy_dq_i_nodelay50;
wire main_nist_clock_ddrphy_dq_i_delayed50;
wire main_nist_clock_ddrphy_dq_t50;
wire main_nist_clock_ddrphy_dq_o_nodelay51;
wire main_nist_clock_ddrphy_dq_o_delayed51;
wire main_nist_clock_ddrphy_dq_i_nodelay51;
wire main_nist_clock_ddrphy_dq_i_delayed51;
wire main_nist_clock_ddrphy_dq_t51;
wire main_nist_clock_ddrphy_dq_o_nodelay52;
wire main_nist_clock_ddrphy_dq_o_delayed52;
wire main_nist_clock_ddrphy_dq_i_nodelay52;
wire main_nist_clock_ddrphy_dq_i_delayed52;
wire main_nist_clock_ddrphy_dq_t52;
wire main_nist_clock_ddrphy_dq_o_nodelay53;
wire main_nist_clock_ddrphy_dq_o_delayed53;
wire main_nist_clock_ddrphy_dq_i_nodelay53;
wire main_nist_clock_ddrphy_dq_i_delayed53;
wire main_nist_clock_ddrphy_dq_t53;
wire main_nist_clock_ddrphy_dq_o_nodelay54;
wire main_nist_clock_ddrphy_dq_o_delayed54;
wire main_nist_clock_ddrphy_dq_i_nodelay54;
wire main_nist_clock_ddrphy_dq_i_delayed54;
wire main_nist_clock_ddrphy_dq_t54;
wire main_nist_clock_ddrphy_dq_o_nodelay55;
wire main_nist_clock_ddrphy_dq_o_delayed55;
wire main_nist_clock_ddrphy_dq_i_nodelay55;
wire main_nist_clock_ddrphy_dq_i_delayed55;
wire main_nist_clock_ddrphy_dq_t55;
wire main_nist_clock_ddrphy_dq_o_nodelay56;
wire main_nist_clock_ddrphy_dq_o_delayed56;
wire main_nist_clock_ddrphy_dq_i_nodelay56;
wire main_nist_clock_ddrphy_dq_i_delayed56;
wire main_nist_clock_ddrphy_dq_t56;
wire main_nist_clock_ddrphy_dq_o_nodelay57;
wire main_nist_clock_ddrphy_dq_o_delayed57;
wire main_nist_clock_ddrphy_dq_i_nodelay57;
wire main_nist_clock_ddrphy_dq_i_delayed57;
wire main_nist_clock_ddrphy_dq_t57;
wire main_nist_clock_ddrphy_dq_o_nodelay58;
wire main_nist_clock_ddrphy_dq_o_delayed58;
wire main_nist_clock_ddrphy_dq_i_nodelay58;
wire main_nist_clock_ddrphy_dq_i_delayed58;
wire main_nist_clock_ddrphy_dq_t58;
wire main_nist_clock_ddrphy_dq_o_nodelay59;
wire main_nist_clock_ddrphy_dq_o_delayed59;
wire main_nist_clock_ddrphy_dq_i_nodelay59;
wire main_nist_clock_ddrphy_dq_i_delayed59;
wire main_nist_clock_ddrphy_dq_t59;
wire main_nist_clock_ddrphy_dq_o_nodelay60;
wire main_nist_clock_ddrphy_dq_o_delayed60;
wire main_nist_clock_ddrphy_dq_i_nodelay60;
wire main_nist_clock_ddrphy_dq_i_delayed60;
wire main_nist_clock_ddrphy_dq_t60;
wire main_nist_clock_ddrphy_dq_o_nodelay61;
wire main_nist_clock_ddrphy_dq_o_delayed61;
wire main_nist_clock_ddrphy_dq_i_nodelay61;
wire main_nist_clock_ddrphy_dq_i_delayed61;
wire main_nist_clock_ddrphy_dq_t61;
wire main_nist_clock_ddrphy_dq_o_nodelay62;
wire main_nist_clock_ddrphy_dq_o_delayed62;
wire main_nist_clock_ddrphy_dq_i_nodelay62;
wire main_nist_clock_ddrphy_dq_i_delayed62;
wire main_nist_clock_ddrphy_dq_t62;
wire main_nist_clock_ddrphy_dq_o_nodelay63;
wire main_nist_clock_ddrphy_dq_o_delayed63;
wire main_nist_clock_ddrphy_dq_i_nodelay63;
wire main_nist_clock_ddrphy_dq_i_delayed63;
wire main_nist_clock_ddrphy_dq_t63;
reg main_nist_clock_ddrphy_n_rddata_en0 = 1'd0;
reg main_nist_clock_ddrphy_n_rddata_en1 = 1'd0;
reg main_nist_clock_ddrphy_n_rddata_en2 = 1'd0;
reg main_nist_clock_ddrphy_n_rddata_en3 = 1'd0;
reg main_nist_clock_ddrphy_n_rddata_en4 = 1'd0;
wire main_nist_clock_ddrphy_oe;
reg [3:0] main_nist_clock_ddrphy_last_wrdata_en = 4'd0;
wire [29:0] main_nist_clock_nist_clock_wb_sdram_adr;
wire [31:0] main_nist_clock_nist_clock_wb_sdram_dat_w;
wire [31:0] main_nist_clock_nist_clock_wb_sdram_dat_r;
wire [3:0] main_nist_clock_nist_clock_wb_sdram_sel;
wire main_nist_clock_nist_clock_wb_sdram_cyc;
wire main_nist_clock_nist_clock_wb_sdram_stb;
wire main_nist_clock_nist_clock_wb_sdram_ack;
wire main_nist_clock_nist_clock_wb_sdram_we;
wire [2:0] main_nist_clock_nist_clock_wb_sdram_cti;
wire [1:0] main_nist_clock_nist_clock_wb_sdram_bte;
wire main_nist_clock_nist_clock_wb_sdram_err;
wire [13:0] main_nist_clock_nist_clock_inti_p0_address;
wire [2:0] main_nist_clock_nist_clock_inti_p0_bank;
reg main_nist_clock_nist_clock_inti_p0_cas_n;
reg main_nist_clock_nist_clock_inti_p0_cs_n;
reg main_nist_clock_nist_clock_inti_p0_ras_n;
reg main_nist_clock_nist_clock_inti_p0_we_n;
wire main_nist_clock_nist_clock_inti_p0_cke;
wire main_nist_clock_nist_clock_inti_p0_odt;
wire main_nist_clock_nist_clock_inti_p0_reset_n;
wire [127:0] main_nist_clock_nist_clock_inti_p0_wrdata;
wire main_nist_clock_nist_clock_inti_p0_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_inti_p0_wrdata_mask;
wire main_nist_clock_nist_clock_inti_p0_rddata_en;
reg [127:0] main_nist_clock_nist_clock_inti_p0_rddata;
reg main_nist_clock_nist_clock_inti_p0_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_inti_p1_address;
wire [2:0] main_nist_clock_nist_clock_inti_p1_bank;
reg main_nist_clock_nist_clock_inti_p1_cas_n;
reg main_nist_clock_nist_clock_inti_p1_cs_n;
reg main_nist_clock_nist_clock_inti_p1_ras_n;
reg main_nist_clock_nist_clock_inti_p1_we_n;
wire main_nist_clock_nist_clock_inti_p1_cke;
wire main_nist_clock_nist_clock_inti_p1_odt;
wire main_nist_clock_nist_clock_inti_p1_reset_n;
wire [127:0] main_nist_clock_nist_clock_inti_p1_wrdata;
wire main_nist_clock_nist_clock_inti_p1_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_inti_p1_wrdata_mask;
wire main_nist_clock_nist_clock_inti_p1_rddata_en;
reg [127:0] main_nist_clock_nist_clock_inti_p1_rddata;
reg main_nist_clock_nist_clock_inti_p1_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_inti_p2_address;
wire [2:0] main_nist_clock_nist_clock_inti_p2_bank;
reg main_nist_clock_nist_clock_inti_p2_cas_n;
reg main_nist_clock_nist_clock_inti_p2_cs_n;
reg main_nist_clock_nist_clock_inti_p2_ras_n;
reg main_nist_clock_nist_clock_inti_p2_we_n;
wire main_nist_clock_nist_clock_inti_p2_cke;
wire main_nist_clock_nist_clock_inti_p2_odt;
wire main_nist_clock_nist_clock_inti_p2_reset_n;
wire [127:0] main_nist_clock_nist_clock_inti_p2_wrdata;
wire main_nist_clock_nist_clock_inti_p2_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_inti_p2_wrdata_mask;
wire main_nist_clock_nist_clock_inti_p2_rddata_en;
reg [127:0] main_nist_clock_nist_clock_inti_p2_rddata;
reg main_nist_clock_nist_clock_inti_p2_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_inti_p3_address;
wire [2:0] main_nist_clock_nist_clock_inti_p3_bank;
reg main_nist_clock_nist_clock_inti_p3_cas_n;
reg main_nist_clock_nist_clock_inti_p3_cs_n;
reg main_nist_clock_nist_clock_inti_p3_ras_n;
reg main_nist_clock_nist_clock_inti_p3_we_n;
wire main_nist_clock_nist_clock_inti_p3_cke;
wire main_nist_clock_nist_clock_inti_p3_odt;
wire main_nist_clock_nist_clock_inti_p3_reset_n;
wire [127:0] main_nist_clock_nist_clock_inti_p3_wrdata;
wire main_nist_clock_nist_clock_inti_p3_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_inti_p3_wrdata_mask;
wire main_nist_clock_nist_clock_inti_p3_rddata_en;
reg [127:0] main_nist_clock_nist_clock_inti_p3_rddata;
reg main_nist_clock_nist_clock_inti_p3_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_slave_p0_address;
wire [2:0] main_nist_clock_nist_clock_slave_p0_bank;
wire main_nist_clock_nist_clock_slave_p0_cas_n;
wire main_nist_clock_nist_clock_slave_p0_cs_n;
wire main_nist_clock_nist_clock_slave_p0_ras_n;
wire main_nist_clock_nist_clock_slave_p0_we_n;
wire main_nist_clock_nist_clock_slave_p0_cke;
wire main_nist_clock_nist_clock_slave_p0_odt;
wire main_nist_clock_nist_clock_slave_p0_reset_n;
wire [127:0] main_nist_clock_nist_clock_slave_p0_wrdata;
wire main_nist_clock_nist_clock_slave_p0_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_slave_p0_wrdata_mask;
wire main_nist_clock_nist_clock_slave_p0_rddata_en;
reg [127:0] main_nist_clock_nist_clock_slave_p0_rddata;
reg main_nist_clock_nist_clock_slave_p0_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_slave_p1_address;
wire [2:0] main_nist_clock_nist_clock_slave_p1_bank;
wire main_nist_clock_nist_clock_slave_p1_cas_n;
wire main_nist_clock_nist_clock_slave_p1_cs_n;
wire main_nist_clock_nist_clock_slave_p1_ras_n;
wire main_nist_clock_nist_clock_slave_p1_we_n;
wire main_nist_clock_nist_clock_slave_p1_cke;
wire main_nist_clock_nist_clock_slave_p1_odt;
wire main_nist_clock_nist_clock_slave_p1_reset_n;
wire [127:0] main_nist_clock_nist_clock_slave_p1_wrdata;
wire main_nist_clock_nist_clock_slave_p1_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_slave_p1_wrdata_mask;
wire main_nist_clock_nist_clock_slave_p1_rddata_en;
reg [127:0] main_nist_clock_nist_clock_slave_p1_rddata;
reg main_nist_clock_nist_clock_slave_p1_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_slave_p2_address;
wire [2:0] main_nist_clock_nist_clock_slave_p2_bank;
wire main_nist_clock_nist_clock_slave_p2_cas_n;
wire main_nist_clock_nist_clock_slave_p2_cs_n;
wire main_nist_clock_nist_clock_slave_p2_ras_n;
wire main_nist_clock_nist_clock_slave_p2_we_n;
wire main_nist_clock_nist_clock_slave_p2_cke;
wire main_nist_clock_nist_clock_slave_p2_odt;
wire main_nist_clock_nist_clock_slave_p2_reset_n;
wire [127:0] main_nist_clock_nist_clock_slave_p2_wrdata;
wire main_nist_clock_nist_clock_slave_p2_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_slave_p2_wrdata_mask;
wire main_nist_clock_nist_clock_slave_p2_rddata_en;
reg [127:0] main_nist_clock_nist_clock_slave_p2_rddata;
reg main_nist_clock_nist_clock_slave_p2_rddata_valid;
wire [13:0] main_nist_clock_nist_clock_slave_p3_address;
wire [2:0] main_nist_clock_nist_clock_slave_p3_bank;
wire main_nist_clock_nist_clock_slave_p3_cas_n;
wire main_nist_clock_nist_clock_slave_p3_cs_n;
wire main_nist_clock_nist_clock_slave_p3_ras_n;
wire main_nist_clock_nist_clock_slave_p3_we_n;
wire main_nist_clock_nist_clock_slave_p3_cke;
wire main_nist_clock_nist_clock_slave_p3_odt;
wire main_nist_clock_nist_clock_slave_p3_reset_n;
wire [127:0] main_nist_clock_nist_clock_slave_p3_wrdata;
wire main_nist_clock_nist_clock_slave_p3_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_slave_p3_wrdata_mask;
wire main_nist_clock_nist_clock_slave_p3_rddata_en;
reg [127:0] main_nist_clock_nist_clock_slave_p3_rddata;
reg main_nist_clock_nist_clock_slave_p3_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_master_p0_address;
reg [2:0] main_nist_clock_nist_clock_master_p0_bank;
reg main_nist_clock_nist_clock_master_p0_cas_n;
reg main_nist_clock_nist_clock_master_p0_cs_n;
reg main_nist_clock_nist_clock_master_p0_ras_n;
reg main_nist_clock_nist_clock_master_p0_we_n;
reg main_nist_clock_nist_clock_master_p0_cke;
reg main_nist_clock_nist_clock_master_p0_odt;
reg main_nist_clock_nist_clock_master_p0_reset_n;
reg [127:0] main_nist_clock_nist_clock_master_p0_wrdata;
reg main_nist_clock_nist_clock_master_p0_wrdata_en;
reg [15:0] main_nist_clock_nist_clock_master_p0_wrdata_mask;
reg main_nist_clock_nist_clock_master_p0_rddata_en;
wire [127:0] main_nist_clock_nist_clock_master_p0_rddata;
wire main_nist_clock_nist_clock_master_p0_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_master_p1_address;
reg [2:0] main_nist_clock_nist_clock_master_p1_bank;
reg main_nist_clock_nist_clock_master_p1_cas_n;
reg main_nist_clock_nist_clock_master_p1_cs_n;
reg main_nist_clock_nist_clock_master_p1_ras_n;
reg main_nist_clock_nist_clock_master_p1_we_n;
reg main_nist_clock_nist_clock_master_p1_cke;
reg main_nist_clock_nist_clock_master_p1_odt;
reg main_nist_clock_nist_clock_master_p1_reset_n;
reg [127:0] main_nist_clock_nist_clock_master_p1_wrdata;
reg main_nist_clock_nist_clock_master_p1_wrdata_en;
reg [15:0] main_nist_clock_nist_clock_master_p1_wrdata_mask;
reg main_nist_clock_nist_clock_master_p1_rddata_en;
wire [127:0] main_nist_clock_nist_clock_master_p1_rddata;
wire main_nist_clock_nist_clock_master_p1_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_master_p2_address;
reg [2:0] main_nist_clock_nist_clock_master_p2_bank;
reg main_nist_clock_nist_clock_master_p2_cas_n;
reg main_nist_clock_nist_clock_master_p2_cs_n;
reg main_nist_clock_nist_clock_master_p2_ras_n;
reg main_nist_clock_nist_clock_master_p2_we_n;
reg main_nist_clock_nist_clock_master_p2_cke;
reg main_nist_clock_nist_clock_master_p2_odt;
reg main_nist_clock_nist_clock_master_p2_reset_n;
reg [127:0] main_nist_clock_nist_clock_master_p2_wrdata;
reg main_nist_clock_nist_clock_master_p2_wrdata_en;
reg [15:0] main_nist_clock_nist_clock_master_p2_wrdata_mask;
reg main_nist_clock_nist_clock_master_p2_rddata_en;
wire [127:0] main_nist_clock_nist_clock_master_p2_rddata;
wire main_nist_clock_nist_clock_master_p2_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_master_p3_address;
reg [2:0] main_nist_clock_nist_clock_master_p3_bank;
reg main_nist_clock_nist_clock_master_p3_cas_n;
reg main_nist_clock_nist_clock_master_p3_cs_n;
reg main_nist_clock_nist_clock_master_p3_ras_n;
reg main_nist_clock_nist_clock_master_p3_we_n;
reg main_nist_clock_nist_clock_master_p3_cke;
reg main_nist_clock_nist_clock_master_p3_odt;
reg main_nist_clock_nist_clock_master_p3_reset_n;
reg [127:0] main_nist_clock_nist_clock_master_p3_wrdata;
reg main_nist_clock_nist_clock_master_p3_wrdata_en;
reg [15:0] main_nist_clock_nist_clock_master_p3_wrdata_mask;
reg main_nist_clock_nist_clock_master_p3_rddata_en;
wire [127:0] main_nist_clock_nist_clock_master_p3_rddata;
wire main_nist_clock_nist_clock_master_p3_rddata_valid;
reg [3:0] main_nist_clock_nist_clock_storage_full = 4'd0;
wire [3:0] main_nist_clock_nist_clock_storage;
reg main_nist_clock_nist_clock_re = 1'd0;
reg [5:0] main_nist_clock_nist_clock_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] main_nist_clock_nist_clock_phaseinjector0_command_storage;
reg main_nist_clock_nist_clock_phaseinjector0_command_re = 1'd0;
wire main_nist_clock_nist_clock_phaseinjector0_command_issue_re;
wire main_nist_clock_nist_clock_phaseinjector0_command_issue_r;
reg main_nist_clock_nist_clock_phaseinjector0_command_issue_w = 1'd0;
reg [13:0] main_nist_clock_nist_clock_phaseinjector0_address_storage_full = 14'd0;
wire [13:0] main_nist_clock_nist_clock_phaseinjector0_address_storage;
reg main_nist_clock_nist_clock_phaseinjector0_address_re = 1'd0;
reg [2:0] main_nist_clock_nist_clock_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] main_nist_clock_nist_clock_phaseinjector0_baddress_storage;
reg main_nist_clock_nist_clock_phaseinjector0_baddress_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full = 128'd0;
wire [127:0] main_nist_clock_nist_clock_phaseinjector0_wrdata_storage;
reg main_nist_clock_nist_clock_phaseinjector0_wrdata_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector0_status = 128'd0;
reg [5:0] main_nist_clock_nist_clock_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] main_nist_clock_nist_clock_phaseinjector1_command_storage;
reg main_nist_clock_nist_clock_phaseinjector1_command_re = 1'd0;
wire main_nist_clock_nist_clock_phaseinjector1_command_issue_re;
wire main_nist_clock_nist_clock_phaseinjector1_command_issue_r;
reg main_nist_clock_nist_clock_phaseinjector1_command_issue_w = 1'd0;
reg [13:0] main_nist_clock_nist_clock_phaseinjector1_address_storage_full = 14'd0;
wire [13:0] main_nist_clock_nist_clock_phaseinjector1_address_storage;
reg main_nist_clock_nist_clock_phaseinjector1_address_re = 1'd0;
reg [2:0] main_nist_clock_nist_clock_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] main_nist_clock_nist_clock_phaseinjector1_baddress_storage;
reg main_nist_clock_nist_clock_phaseinjector1_baddress_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full = 128'd0;
wire [127:0] main_nist_clock_nist_clock_phaseinjector1_wrdata_storage;
reg main_nist_clock_nist_clock_phaseinjector1_wrdata_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector1_status = 128'd0;
reg [5:0] main_nist_clock_nist_clock_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] main_nist_clock_nist_clock_phaseinjector2_command_storage;
reg main_nist_clock_nist_clock_phaseinjector2_command_re = 1'd0;
wire main_nist_clock_nist_clock_phaseinjector2_command_issue_re;
wire main_nist_clock_nist_clock_phaseinjector2_command_issue_r;
reg main_nist_clock_nist_clock_phaseinjector2_command_issue_w = 1'd0;
reg [13:0] main_nist_clock_nist_clock_phaseinjector2_address_storage_full = 14'd0;
wire [13:0] main_nist_clock_nist_clock_phaseinjector2_address_storage;
reg main_nist_clock_nist_clock_phaseinjector2_address_re = 1'd0;
reg [2:0] main_nist_clock_nist_clock_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] main_nist_clock_nist_clock_phaseinjector2_baddress_storage;
reg main_nist_clock_nist_clock_phaseinjector2_baddress_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full = 128'd0;
wire [127:0] main_nist_clock_nist_clock_phaseinjector2_wrdata_storage;
reg main_nist_clock_nist_clock_phaseinjector2_wrdata_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector2_status = 128'd0;
reg [5:0] main_nist_clock_nist_clock_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] main_nist_clock_nist_clock_phaseinjector3_command_storage;
reg main_nist_clock_nist_clock_phaseinjector3_command_re = 1'd0;
wire main_nist_clock_nist_clock_phaseinjector3_command_issue_re;
wire main_nist_clock_nist_clock_phaseinjector3_command_issue_r;
reg main_nist_clock_nist_clock_phaseinjector3_command_issue_w = 1'd0;
reg [13:0] main_nist_clock_nist_clock_phaseinjector3_address_storage_full = 14'd0;
wire [13:0] main_nist_clock_nist_clock_phaseinjector3_address_storage;
reg main_nist_clock_nist_clock_phaseinjector3_address_re = 1'd0;
reg [2:0] main_nist_clock_nist_clock_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] main_nist_clock_nist_clock_phaseinjector3_baddress_storage;
reg main_nist_clock_nist_clock_phaseinjector3_baddress_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full = 128'd0;
wire [127:0] main_nist_clock_nist_clock_phaseinjector3_wrdata_storage;
reg main_nist_clock_nist_clock_phaseinjector3_wrdata_re = 1'd0;
reg [127:0] main_nist_clock_nist_clock_phaseinjector3_status = 128'd0;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_dfi_p0_address;
wire [2:0] main_nist_clock_nist_clock_sdram_controller_dfi_p0_bank;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p0_cs_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p0_cke;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p0_odt;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p0_reset_n;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata_en = 1'd0;
wire [15:0] main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata_mask;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_en;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_dfi_p1_address;
wire [2:0] main_nist_clock_nist_clock_sdram_controller_dfi_p1_bank;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p1_cas_n = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p1_cs_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p1_ras_n = 1'd1;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p1_we_n = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p1_cke;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p1_odt;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p1_reset_n;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata_en = 1'd0;
wire [15:0] main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata_mask;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata_en = 1'd0;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_dfi_p2_address;
wire [2:0] main_nist_clock_nist_clock_sdram_controller_dfi_p2_bank;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p2_cas_n;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p2_cs_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p2_ras_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p2_we_n;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p2_cke;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p2_odt;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p2_reset_n;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_en;
wire [15:0] main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_mask;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata_en = 1'd0;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata_valid;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_dfi_p3_address;
wire [2:0] main_nist_clock_nist_clock_sdram_controller_dfi_p3_bank;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p3_cas_n = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p3_cs_n;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p3_ras_n = 1'd1;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p3_we_n = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p3_cke;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p3_odt;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p3_reset_n;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata_en = 1'd0;
wire [15:0] main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata_mask;
reg main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata_en = 1'd0;
wire [127:0] main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata;
wire main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata_valid;
wire [29:0] main_nist_clock_nist_clock_sdram_controller_bus_adr;
wire [511:0] main_nist_clock_nist_clock_sdram_controller_bus_dat_w;
wire [511:0] main_nist_clock_nist_clock_sdram_controller_bus_dat_r;
wire [63:0] main_nist_clock_nist_clock_sdram_controller_bus_sel;
wire main_nist_clock_nist_clock_sdram_controller_bus_cyc;
wire main_nist_clock_nist_clock_sdram_controller_bus_stb;
reg main_nist_clock_nist_clock_sdram_controller_bus_ack;
wire main_nist_clock_nist_clock_sdram_controller_bus_we;
wire [2:0] main_nist_clock_nist_clock_sdram_controller_bus_cti;
wire [1:0] main_nist_clock_nist_clock_sdram_controller_bus_bte;
reg main_nist_clock_nist_clock_sdram_controller_bus_err = 1'd0;
reg main_nist_clock_nist_clock_sdram_controller_precharge_all;
reg main_nist_clock_nist_clock_sdram_controller_activate;
reg main_nist_clock_nist_clock_sdram_controller_refresh;
reg main_nist_clock_nist_clock_sdram_controller_write;
reg main_nist_clock_nist_clock_sdram_controller_read;
wire main_nist_clock_nist_clock_sdram_controller_bank_idle;
wire main_nist_clock_nist_clock_sdram_controller_bank_hit;
wire main_nist_clock_nist_clock_sdram_controller_bank0_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank0_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank0_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank0_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank0_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce0;
wire main_nist_clock_nist_clock_sdram_controller_reset0;
wire main_nist_clock_nist_clock_sdram_controller_bank1_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank1_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank1_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank1_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank1_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce1;
wire main_nist_clock_nist_clock_sdram_controller_reset1;
wire main_nist_clock_nist_clock_sdram_controller_bank2_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank2_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank2_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank2_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank2_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce2;
wire main_nist_clock_nist_clock_sdram_controller_reset2;
wire main_nist_clock_nist_clock_sdram_controller_bank3_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank3_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank3_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank3_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank3_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce3;
wire main_nist_clock_nist_clock_sdram_controller_reset3;
wire main_nist_clock_nist_clock_sdram_controller_bank4_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank4_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank4_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank4_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank4_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce4;
wire main_nist_clock_nist_clock_sdram_controller_reset4;
wire main_nist_clock_nist_clock_sdram_controller_bank5_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank5_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank5_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank5_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank5_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce5;
wire main_nist_clock_nist_clock_sdram_controller_reset5;
wire main_nist_clock_nist_clock_sdram_controller_bank6_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank6_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank6_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank6_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank6_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce6;
wire main_nist_clock_nist_clock_sdram_controller_reset6;
wire main_nist_clock_nist_clock_sdram_controller_bank7_open;
wire [13:0] main_nist_clock_nist_clock_sdram_controller_bank7_row0;
reg main_nist_clock_nist_clock_sdram_controller_bank7_idle = 1'd1;
wire main_nist_clock_nist_clock_sdram_controller_bank7_hit;
reg [13:0] main_nist_clock_nist_clock_sdram_controller_bank7_row1 = 14'd0;
reg main_nist_clock_nist_clock_sdram_controller_ce7;
wire main_nist_clock_nist_clock_sdram_controller_reset7;
wire main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_wait;
wire main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_done;
reg [2:0] main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count = 3'd4;
wire main_nist_clock_nist_clock_sdram_controller_refresh_timer_wait;
wire main_nist_clock_nist_clock_sdram_controller_refresh_timer_done;
reg [9:0] main_nist_clock_nist_clock_sdram_controller_refresh_timer_count = 10'd975;
wire [29:0] main_nist_clock_nist_clock_bridge_if_bus_adr;
wire [511:0] main_nist_clock_nist_clock_bridge_if_bus_dat_w;
wire [511:0] main_nist_clock_nist_clock_bridge_if_bus_dat_r;
wire [63:0] main_nist_clock_nist_clock_bridge_if_bus_sel;
reg main_nist_clock_nist_clock_bridge_if_bus_cyc;
reg main_nist_clock_nist_clock_bridge_if_bus_stb;
wire main_nist_clock_nist_clock_bridge_if_bus_ack;
reg main_nist_clock_nist_clock_bridge_if_bus_we;
reg [2:0] main_nist_clock_nist_clock_bridge_if_bus_cti = 3'd0;
reg [1:0] main_nist_clock_nist_clock_bridge_if_bus_bte = 2'd0;
wire main_nist_clock_nist_clock_bridge_if_bus_err;
wire [10:0] main_nist_clock_nist_clock_data_port_adr;
wire [511:0] main_nist_clock_nist_clock_data_port_dat_r;
reg [63:0] main_nist_clock_nist_clock_data_port_we;
reg [511:0] main_nist_clock_nist_clock_data_port_dat_w;
reg main_nist_clock_nist_clock_write_from_slave;
reg [3:0] main_nist_clock_nist_clock_adr_offset_r = 4'd0;
wire [10:0] main_nist_clock_nist_clock_tag_port_adr;
wire [23:0] main_nist_clock_nist_clock_tag_port_dat_r;
reg main_nist_clock_nist_clock_tag_port_we;
wire [23:0] main_nist_clock_nist_clock_tag_port_dat_w;
wire [22:0] main_nist_clock_nist_clock_tag_do_tag;
wire main_nist_clock_nist_clock_tag_do_dirty;
wire [22:0] main_nist_clock_nist_clock_tag_di_tag;
reg main_nist_clock_nist_clock_tag_di_dirty;
reg main_nist_clock_nist_clock_word_clr;
reg main_nist_clock_nist_clock_word_inc;
reg main_nist_clock_clk;
wire [29:0] main_nist_clock_spiflash_bus_adr;
wire [31:0] main_nist_clock_spiflash_bus_dat_w;
wire [31:0] main_nist_clock_spiflash_bus_dat_r;
wire [3:0] main_nist_clock_spiflash_bus_sel;
wire main_nist_clock_spiflash_bus_cyc;
wire main_nist_clock_spiflash_bus_stb;
reg main_nist_clock_spiflash_bus_ack = 1'd0;
wire main_nist_clock_spiflash_bus_we;
wire [2:0] main_nist_clock_spiflash_bus_cti;
wire [1:0] main_nist_clock_spiflash_bus_bte;
reg main_nist_clock_spiflash_bus_err = 1'd0;
reg [3:0] main_nist_clock_spiflash_bitbang_storage_full = 4'd0;
wire [3:0] main_nist_clock_spiflash_bitbang_storage;
reg main_nist_clock_spiflash_bitbang_re = 1'd0;
reg main_nist_clock_spiflash_status;
reg main_nist_clock_spiflash_bitbang_en_storage_full = 1'd0;
wire main_nist_clock_spiflash_bitbang_en_storage;
reg main_nist_clock_spiflash_bitbang_en_re = 1'd0;
reg main_nist_clock_spiflash_cs_n1 = 1'd1;
reg main_nist_clock_spiflash_clk = 1'd0;
reg main_nist_clock_spiflash_dq_oe = 1'd0;
reg [3:0] main_nist_clock_spiflash_o;
reg main_nist_clock_spiflash_oe;
wire [3:0] main_nist_clock_spiflash_i0;
reg [31:0] main_nist_clock_spiflash_sr = 32'd0;
reg main_nist_clock_spiflash_i1 = 1'd0;
reg [3:0] main_nist_clock_spiflash_dqi = 4'd0;
reg [6:0] main_nist_clock_spiflash_counter = 7'd0;
reg main_ethphy_mode0 = 1'd0;
wire main_ethphy_mode_status;
reg main_ethphy_mode1;
reg main_ethphy_update_mode;
wire main_ethphy_eth_tick;
reg [9:0] main_ethphy_eth_counter = 10'd0;
wire main_ethphy_sys_tick;
wire main_ethphy_i;
wire main_ethphy_o;
reg main_ethphy_toggle_i = 1'd0;
wire main_ethphy_toggle_o;
reg main_ethphy_toggle_o_r = 1'd0;
reg [23:0] main_ethphy_sys_counter = 24'd0;
reg main_ethphy_sys_counter_reset;
reg main_ethphy_sys_counter_ce;
reg main_ethphy_storage_full = 1'd0;
wire main_ethphy_storage;
reg main_ethphy_re = 1'd0;
wire eth_rx_clk;
wire eth_rx_rst;
wire eth_tx_clk;
wire eth_tx_rst;
wire main_ethphy_liteethphygmiimiitx_sink_sink_stb0;
wire main_ethphy_liteethphygmiimiitx_sink_sink_ack0;
wire main_ethphy_liteethphygmiimiitx_sink_sink_eop0;
wire [7:0] main_ethphy_liteethphygmiimiitx_sink_sink_payload_data0;
wire main_ethphy_liteethphygmiimiitx_sink_sink_payload_last_be0;
wire main_ethphy_liteethphygmiimiitx_sink_sink_payload_error0;
reg main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_er = 1'd0;
reg main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_en = 1'd0;
reg [7:0] main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_data = 8'd0;
wire main_ethphy_liteethphygmiimiitx_gmii_tx_sink_stb;
reg main_ethphy_liteethphygmiimiitx_gmii_tx_sink_ack = 1'd0;
wire main_ethphy_liteethphygmiimiitx_gmii_tx_sink_eop;
wire [7:0] main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_data;
wire main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_last_be;
wire main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_error;
reg main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_er = 1'd0;
reg main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_en = 1'd0;
reg [7:0] main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_data = 8'd0;
wire main_ethphy_liteethphygmiimiitx_sink_sink_stb1;
wire main_ethphy_liteethphygmiimiitx_sink_sink_ack1;
wire main_ethphy_liteethphygmiimiitx_sink_sink_eop1;
wire [7:0] main_ethphy_liteethphygmiimiitx_sink_sink_payload_data1;
wire main_ethphy_liteethphygmiimiitx_sink_sink_payload_last_be1;
wire main_ethphy_liteethphygmiimiitx_sink_sink_payload_error1;
wire main_ethphy_liteethphygmiimiitx_converter_sink_stb;
wire main_ethphy_liteethphygmiimiitx_converter_sink_ack;
reg main_ethphy_liteethphygmiimiitx_converter_sink_eop = 1'd0;
wire [7:0] main_ethphy_liteethphygmiimiitx_converter_sink_payload_data;
wire main_ethphy_liteethphygmiimiitx_converter_source_stb;
wire main_ethphy_liteethphygmiimiitx_converter_source_ack;
wire main_ethphy_liteethphygmiimiitx_converter_source_eop;
reg [3:0] main_ethphy_liteethphygmiimiitx_converter_source_payload_data;
reg main_ethphy_liteethphygmiimiitx_converter_mux = 1'd0;
wire main_ethphy_liteethphygmiimiitx_converter_last;
wire main_ethphy_liteethphygmiimiitx_demux_sink_stb;
reg main_ethphy_liteethphygmiimiitx_demux_sink_ack;
wire main_ethphy_liteethphygmiimiitx_demux_sink_eop;
wire [7:0] main_ethphy_liteethphygmiimiitx_demux_sink_payload_data;
wire main_ethphy_liteethphygmiimiitx_demux_sink_payload_last_be;
wire main_ethphy_liteethphygmiimiitx_demux_sink_payload_error;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_stb;
wire main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_ack;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_eop;
reg [7:0] main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_data;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_last_be;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_error;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_stb;
wire main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_ack;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_eop;
reg [7:0] main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_data;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_last_be;
reg main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_error;
wire main_ethphy_liteethphygmiimiitx_demux_sel;
wire main_ethphy_liteethphygmiimiirx_source_source_stb0;
wire main_ethphy_liteethphygmiimiirx_source_source_ack0;
wire main_ethphy_liteethphygmiimiirx_source_source_eop0;
wire [7:0] main_ethphy_liteethphygmiimiirx_source_source_payload_data0;
wire main_ethphy_liteethphygmiimiirx_source_source_payload_last_be0;
wire main_ethphy_liteethphygmiimiirx_source_source_payload_error0;
reg main_ethphy_liteethphygmiimiirx_pads_d_rx_dv = 1'd0;
reg [7:0] main_ethphy_liteethphygmiimiirx_pads_d_rx_data = 8'd0;
reg main_ethphy_liteethphygmiimiirx_gmii_rx_source_stb = 1'd0;
wire main_ethphy_liteethphygmiimiirx_gmii_rx_source_ack;
wire main_ethphy_liteethphygmiimiirx_gmii_rx_source_eop;
reg [7:0] main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_data = 8'd0;
reg main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_last_be = 1'd0;
reg main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_error = 1'd0;
reg main_ethphy_liteethphygmiimiirx_gmii_rx_rx_dv_d = 1'd0;
wire main_ethphy_liteethphygmiimiirx_source_source_stb1;
wire main_ethphy_liteethphygmiimiirx_source_source_ack1;
wire main_ethphy_liteethphygmiimiirx_source_source_eop1;
wire [7:0] main_ethphy_liteethphygmiimiirx_source_source_payload_data1;
reg main_ethphy_liteethphygmiimiirx_source_source_payload_last_be1 = 1'd0;
reg main_ethphy_liteethphygmiimiirx_source_source_payload_error1 = 1'd0;
reg main_ethphy_liteethphygmiimiirx_converter_sink_stb = 1'd0;
wire main_ethphy_liteethphygmiimiirx_converter_sink_ack;
wire main_ethphy_liteethphygmiimiirx_converter_sink_eop;
reg [3:0] main_ethphy_liteethphygmiimiirx_converter_sink_payload_data = 4'd0;
wire main_ethphy_liteethphygmiimiirx_converter_source_stb;
wire main_ethphy_liteethphygmiimiirx_converter_source_ack;
reg main_ethphy_liteethphygmiimiirx_converter_source_eop = 1'd0;
reg [7:0] main_ethphy_liteethphygmiimiirx_converter_source_payload_data = 8'd0;
reg main_ethphy_liteethphygmiimiirx_converter_demux = 1'd0;
wire main_ethphy_liteethphygmiimiirx_converter_load_part;
reg main_ethphy_liteethphygmiimiirx_converter_strobe_all = 1'd0;
reg main_ethphy_liteethphygmiimiirx_converter_reset = 1'd0;
reg main_ethphy_liteethphygmiimiirx_mux_source_stb;
wire main_ethphy_liteethphygmiimiirx_mux_source_ack;
reg main_ethphy_liteethphygmiimiirx_mux_source_eop;
reg [7:0] main_ethphy_liteethphygmiimiirx_mux_source_payload_data;
reg main_ethphy_liteethphygmiimiirx_mux_source_payload_last_be;
reg main_ethphy_liteethphygmiimiirx_mux_source_payload_error;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_stb;
reg main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_ack;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_eop;
wire [7:0] main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_data;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_last_be;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_error;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_stb;
reg main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_ack;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_eop;
wire [7:0] main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_data;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_last_be;
wire main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_error;
wire main_ethphy_liteethphygmiimiirx_mux_sel;
wire main_tx_gap_inserter_sink_stb;
reg main_tx_gap_inserter_sink_ack;
wire main_tx_gap_inserter_sink_eop;
wire [7:0] main_tx_gap_inserter_sink_payload_data;
wire main_tx_gap_inserter_sink_payload_last_be;
wire main_tx_gap_inserter_sink_payload_error;
reg main_tx_gap_inserter_source_stb;
wire main_tx_gap_inserter_source_ack;
reg main_tx_gap_inserter_source_eop;
reg [7:0] main_tx_gap_inserter_source_payload_data;
reg main_tx_gap_inserter_source_payload_last_be;
reg main_tx_gap_inserter_source_payload_error;
reg [3:0] main_tx_gap_inserter_counter = 4'd0;
reg main_tx_gap_inserter_counter_reset;
reg main_tx_gap_inserter_counter_ce;
reg [31:0] main_preamble_errors_status = 32'd0;
reg [31:0] main_crc_errors_status = 32'd0;
wire main_preamble_inserter_sink_stb;
reg main_preamble_inserter_sink_ack;
wire main_preamble_inserter_sink_eop;
wire [7:0] main_preamble_inserter_sink_payload_data;
wire main_preamble_inserter_sink_payload_last_be;
wire main_preamble_inserter_sink_payload_error;
reg main_preamble_inserter_source_stb;
wire main_preamble_inserter_source_ack;
reg main_preamble_inserter_source_eop;
reg [7:0] main_preamble_inserter_source_payload_data;
wire main_preamble_inserter_source_payload_last_be;
reg main_preamble_inserter_source_payload_error;
reg [63:0] main_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] main_preamble_inserter_cnt = 3'd0;
reg main_preamble_inserter_clr_cnt;
reg main_preamble_inserter_inc_cnt;
wire main_preamble_checker_sink_stb;
reg main_preamble_checker_sink_ack;
wire main_preamble_checker_sink_eop;
wire [7:0] main_preamble_checker_sink_payload_data;
wire main_preamble_checker_sink_payload_last_be;
wire main_preamble_checker_sink_payload_error;
reg main_preamble_checker_source_stb;
wire main_preamble_checker_source_ack;
reg main_preamble_checker_source_eop;
wire [7:0] main_preamble_checker_source_payload_data;
wire main_preamble_checker_source_payload_last_be;
reg main_preamble_checker_source_payload_error;
reg main_preamble_checker_error;
wire main_crc32_inserter_sink_stb;
reg main_crc32_inserter_sink_ack;
wire main_crc32_inserter_sink_eop;
wire [7:0] main_crc32_inserter_sink_payload_data;
wire main_crc32_inserter_sink_payload_last_be;
wire main_crc32_inserter_sink_payload_error;
reg main_crc32_inserter_source_stb;
wire main_crc32_inserter_source_ack;
reg main_crc32_inserter_source_eop;
reg [7:0] main_crc32_inserter_source_payload_data;
reg main_crc32_inserter_source_payload_last_be;
reg main_crc32_inserter_source_payload_error;
reg [7:0] main_crc32_inserter_data0;
wire [31:0] main_crc32_inserter_value;
wire main_crc32_inserter_error;
wire [7:0] main_crc32_inserter_data1;
wire [31:0] main_crc32_inserter_last;
reg [31:0] main_crc32_inserter_next;
reg [31:0] main_crc32_inserter_reg = 32'd4294967295;
reg main_crc32_inserter_ce;
reg main_crc32_inserter_reset;
reg [1:0] main_crc32_inserter_cnt = 2'd3;
wire main_crc32_inserter_cnt_done;
reg main_crc32_inserter_is_ongoing0;
reg main_crc32_inserter_is_ongoing1;
wire main_crc32_checker_sink_sink_stb;
reg main_crc32_checker_sink_sink_ack;
wire main_crc32_checker_sink_sink_eop;
wire [7:0] main_crc32_checker_sink_sink_payload_data;
wire main_crc32_checker_sink_sink_payload_last_be;
wire main_crc32_checker_sink_sink_payload_error;
wire main_crc32_checker_source_source_stb;
wire main_crc32_checker_source_source_ack;
wire main_crc32_checker_source_source_eop;
wire [7:0] main_crc32_checker_source_source_payload_data;
wire main_crc32_checker_source_source_payload_last_be;
reg main_crc32_checker_source_source_payload_error;
wire main_crc32_checker_error;
wire [7:0] main_crc32_checker_crc_data0;
wire [31:0] main_crc32_checker_crc_value;
wire main_crc32_checker_crc_error;
wire [7:0] main_crc32_checker_crc_data1;
wire [31:0] main_crc32_checker_crc_last;
reg [31:0] main_crc32_checker_crc_next;
reg [31:0] main_crc32_checker_crc_reg = 32'd4294967295;
reg main_crc32_checker_crc_ce;
reg main_crc32_checker_crc_reset;
reg main_crc32_checker_syncfifo_sink_stb;
wire main_crc32_checker_syncfifo_sink_ack;
wire main_crc32_checker_syncfifo_sink_eop;
wire [7:0] main_crc32_checker_syncfifo_sink_payload_data;
wire main_crc32_checker_syncfifo_sink_payload_last_be;
wire main_crc32_checker_syncfifo_sink_payload_error;
wire main_crc32_checker_syncfifo_source_stb;
wire main_crc32_checker_syncfifo_source_ack;
wire main_crc32_checker_syncfifo_source_eop;
wire [7:0] main_crc32_checker_syncfifo_source_payload_data;
wire main_crc32_checker_syncfifo_source_payload_last_be;
wire main_crc32_checker_syncfifo_source_payload_error;
wire main_crc32_checker_syncfifo_syncfifo_we;
wire main_crc32_checker_syncfifo_syncfifo_writable;
wire main_crc32_checker_syncfifo_syncfifo_re;
wire main_crc32_checker_syncfifo_syncfifo_readable;
wire [10:0] main_crc32_checker_syncfifo_syncfifo_din;
wire [10:0] main_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] main_crc32_checker_syncfifo_level = 3'd0;
reg main_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] main_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] main_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] main_crc32_checker_syncfifo_wrport_adr;
wire [10:0] main_crc32_checker_syncfifo_wrport_dat_r;
wire main_crc32_checker_syncfifo_wrport_we;
wire [10:0] main_crc32_checker_syncfifo_wrport_dat_w;
wire main_crc32_checker_syncfifo_do_read;
wire [2:0] main_crc32_checker_syncfifo_rdport_adr;
wire [10:0] main_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] main_crc32_checker_syncfifo_fifo_in_payload_data;
wire main_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire main_crc32_checker_syncfifo_fifo_in_payload_error;
wire main_crc32_checker_syncfifo_fifo_in_eop;
wire [7:0] main_crc32_checker_syncfifo_fifo_out_payload_data;
wire main_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire main_crc32_checker_syncfifo_fifo_out_payload_error;
wire main_crc32_checker_syncfifo_fifo_out_eop;
reg main_crc32_checker_fifo_reset;
wire main_crc32_checker_fifo_in;
wire main_crc32_checker_fifo_out;
wire main_crc32_checker_fifo_full;
wire main_ps_preamble_error_i;
wire main_ps_preamble_error_o;
reg main_ps_preamble_error_toggle_i = 1'd0;
wire main_ps_preamble_error_toggle_o;
reg main_ps_preamble_error_toggle_o_r = 1'd0;
wire main_ps_crc_error_i;
wire main_ps_crc_error_o;
reg main_ps_crc_error_toggle_i = 1'd0;
wire main_ps_crc_error_toggle_o;
reg main_ps_crc_error_toggle_o_r = 1'd0;
wire main_padding_inserter_sink_stb;
reg main_padding_inserter_sink_ack;
wire main_padding_inserter_sink_eop;
wire [7:0] main_padding_inserter_sink_payload_data;
wire main_padding_inserter_sink_payload_last_be;
wire main_padding_inserter_sink_payload_error;
reg main_padding_inserter_source_stb;
wire main_padding_inserter_source_ack;
reg main_padding_inserter_source_eop;
reg [7:0] main_padding_inserter_source_payload_data;
reg main_padding_inserter_source_payload_last_be;
reg main_padding_inserter_source_payload_error;
reg [15:0] main_padding_inserter_counter = 16'd1;
wire main_padding_inserter_counter_done;
reg main_padding_inserter_counter_reset;
reg main_padding_inserter_counter_ce;
wire main_padding_checker_sink_stb;
wire main_padding_checker_sink_ack;
wire main_padding_checker_sink_eop;
wire [7:0] main_padding_checker_sink_payload_data;
wire main_padding_checker_sink_payload_last_be;
wire main_padding_checker_sink_payload_error;
wire main_padding_checker_source_stb;
wire main_padding_checker_source_ack;
wire main_padding_checker_source_eop;
wire [7:0] main_padding_checker_source_payload_data;
wire main_padding_checker_source_payload_last_be;
wire main_padding_checker_source_payload_error;
wire main_tx_last_be_sink_stb;
wire main_tx_last_be_sink_ack;
wire main_tx_last_be_sink_eop;
wire [7:0] main_tx_last_be_sink_payload_data;
wire main_tx_last_be_sink_payload_last_be;
wire main_tx_last_be_sink_payload_error;
wire main_tx_last_be_source_stb;
wire main_tx_last_be_source_ack;
wire main_tx_last_be_source_eop;
wire [7:0] main_tx_last_be_source_payload_data;
reg main_tx_last_be_source_payload_last_be = 1'd0;
reg main_tx_last_be_source_payload_error = 1'd0;
reg main_tx_last_be_ongoing = 1'd1;
wire main_rx_last_be_sink_stb;
wire main_rx_last_be_sink_ack;
wire main_rx_last_be_sink_eop;
wire [7:0] main_rx_last_be_sink_payload_data;
wire main_rx_last_be_sink_payload_last_be;
wire main_rx_last_be_sink_payload_error;
wire main_rx_last_be_source_stb;
wire main_rx_last_be_source_ack;
wire main_rx_last_be_source_eop;
wire [7:0] main_rx_last_be_source_payload_data;
reg main_rx_last_be_source_payload_last_be;
wire main_rx_last_be_source_payload_error;
wire main_tx_converter_sink_sink_stb;
wire main_tx_converter_sink_sink_ack;
wire main_tx_converter_sink_sink_eop;
wire [31:0] main_tx_converter_sink_sink_payload_data;
wire [3:0] main_tx_converter_sink_sink_payload_last_be;
wire [3:0] main_tx_converter_sink_sink_payload_error;
wire main_tx_converter_source_source_stb;
wire main_tx_converter_source_source_ack;
wire main_tx_converter_source_source_eop;
wire [7:0] main_tx_converter_source_source_payload_data;
wire main_tx_converter_source_source_payload_last_be;
wire main_tx_converter_source_source_payload_error;
wire main_tx_converter_converter_sink_stb;
wire main_tx_converter_converter_sink_ack;
wire main_tx_converter_converter_sink_eop;
reg [39:0] main_tx_converter_converter_sink_payload_data;
wire main_tx_converter_converter_source_stb;
wire main_tx_converter_converter_source_ack;
wire main_tx_converter_converter_source_eop;
reg [9:0] main_tx_converter_converter_source_payload_data;
reg [1:0] main_tx_converter_converter_mux = 2'd0;
wire main_tx_converter_converter_last;
wire main_rx_converter_sink_sink_stb;
wire main_rx_converter_sink_sink_ack;
wire main_rx_converter_sink_sink_eop;
wire [7:0] main_rx_converter_sink_sink_payload_data;
wire main_rx_converter_sink_sink_payload_last_be;
wire main_rx_converter_sink_sink_payload_error;
wire main_rx_converter_source_source_stb;
wire main_rx_converter_source_source_ack;
wire main_rx_converter_source_source_eop;
reg [31:0] main_rx_converter_source_source_payload_data;
reg [3:0] main_rx_converter_source_source_payload_last_be;
reg [3:0] main_rx_converter_source_source_payload_error;
wire main_rx_converter_converter_sink_stb;
wire main_rx_converter_converter_sink_ack;
wire main_rx_converter_converter_sink_eop;
wire [9:0] main_rx_converter_converter_sink_payload_data;
wire main_rx_converter_converter_source_stb;
wire main_rx_converter_converter_source_ack;
reg main_rx_converter_converter_source_eop = 1'd0;
reg [39:0] main_rx_converter_converter_source_payload_data = 40'd0;
reg [1:0] main_rx_converter_converter_demux = 2'd0;
wire main_rx_converter_converter_load_part;
reg main_rx_converter_converter_strobe_all = 1'd0;
wire main_tx_cdc_sink_stb;
wire main_tx_cdc_sink_ack;
wire main_tx_cdc_sink_eop;
wire [31:0] main_tx_cdc_sink_payload_data;
wire [3:0] main_tx_cdc_sink_payload_last_be;
wire [3:0] main_tx_cdc_sink_payload_error;
wire main_tx_cdc_source_stb;
wire main_tx_cdc_source_ack;
wire main_tx_cdc_source_eop;
wire [31:0] main_tx_cdc_source_payload_data;
wire [3:0] main_tx_cdc_source_payload_last_be;
wire [3:0] main_tx_cdc_source_payload_error;
wire main_tx_cdc_asyncfifo_we;
wire main_tx_cdc_asyncfifo_writable;
wire main_tx_cdc_asyncfifo_re;
wire main_tx_cdc_asyncfifo_readable;
wire [40:0] main_tx_cdc_asyncfifo_din;
wire [40:0] main_tx_cdc_asyncfifo_dout;
wire main_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_tx_cdc_graycounter0_q_next;
reg [6:0] main_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_tx_cdc_graycounter0_q_next_binary;
wire main_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_tx_cdc_graycounter1_q_next;
reg [6:0] main_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_tx_cdc_graycounter1_q_next_binary;
wire [6:0] main_tx_cdc_produce_rdomain;
wire [6:0] main_tx_cdc_consume_wdomain;
wire [5:0] main_tx_cdc_wrport_adr;
wire [40:0] main_tx_cdc_wrport_dat_r;
wire main_tx_cdc_wrport_we;
wire [40:0] main_tx_cdc_wrport_dat_w;
wire [5:0] main_tx_cdc_rdport_adr;
wire [40:0] main_tx_cdc_rdport_dat_r;
wire [31:0] main_tx_cdc_fifo_in_payload_data;
wire [3:0] main_tx_cdc_fifo_in_payload_last_be;
wire [3:0] main_tx_cdc_fifo_in_payload_error;
wire main_tx_cdc_fifo_in_eop;
wire [31:0] main_tx_cdc_fifo_out_payload_data;
wire [3:0] main_tx_cdc_fifo_out_payload_last_be;
wire [3:0] main_tx_cdc_fifo_out_payload_error;
wire main_tx_cdc_fifo_out_eop;
wire main_rx_cdc_sink_stb;
wire main_rx_cdc_sink_ack;
wire main_rx_cdc_sink_eop;
wire [31:0] main_rx_cdc_sink_payload_data;
wire [3:0] main_rx_cdc_sink_payload_last_be;
wire [3:0] main_rx_cdc_sink_payload_error;
wire main_rx_cdc_source_stb;
wire main_rx_cdc_source_ack;
wire main_rx_cdc_source_eop;
wire [31:0] main_rx_cdc_source_payload_data;
wire [3:0] main_rx_cdc_source_payload_last_be;
wire [3:0] main_rx_cdc_source_payload_error;
wire main_rx_cdc_asyncfifo_we;
wire main_rx_cdc_asyncfifo_writable;
wire main_rx_cdc_asyncfifo_re;
wire main_rx_cdc_asyncfifo_readable;
wire [40:0] main_rx_cdc_asyncfifo_din;
wire [40:0] main_rx_cdc_asyncfifo_dout;
wire main_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] main_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] main_rx_cdc_graycounter0_q_next;
reg [6:0] main_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] main_rx_cdc_graycounter0_q_next_binary;
wire main_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] main_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] main_rx_cdc_graycounter1_q_next;
reg [6:0] main_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] main_rx_cdc_graycounter1_q_next_binary;
wire [6:0] main_rx_cdc_produce_rdomain;
wire [6:0] main_rx_cdc_consume_wdomain;
wire [5:0] main_rx_cdc_wrport_adr;
wire [40:0] main_rx_cdc_wrport_dat_r;
wire main_rx_cdc_wrport_we;
wire [40:0] main_rx_cdc_wrport_dat_w;
wire [5:0] main_rx_cdc_rdport_adr;
wire [40:0] main_rx_cdc_rdport_dat_r;
wire [31:0] main_rx_cdc_fifo_in_payload_data;
wire [3:0] main_rx_cdc_fifo_in_payload_last_be;
wire [3:0] main_rx_cdc_fifo_in_payload_error;
wire main_rx_cdc_fifo_in_eop;
wire [31:0] main_rx_cdc_fifo_out_payload_data;
wire [3:0] main_rx_cdc_fifo_out_payload_last_be;
wire [3:0] main_rx_cdc_fifo_out_payload_error;
wire main_rx_cdc_fifo_out_eop;
wire main_sink_stb;
wire main_sink_ack;
wire main_sink_eop;
wire [31:0] main_sink_payload_data;
wire [3:0] main_sink_payload_last_be;
wire [3:0] main_sink_payload_error;
wire main_source_stb;
wire main_source_ack;
wire main_source_eop;
wire [31:0] main_source_payload_data;
wire [3:0] main_source_payload_last_be;
wire [3:0] main_source_payload_error;
wire [29:0] main_bus_adr;
wire [31:0] main_bus_dat_w;
wire [31:0] main_bus_dat_r;
wire [3:0] main_bus_sel;
wire main_bus_cyc;
wire main_bus_stb;
wire main_bus_ack;
wire main_bus_we;
wire [2:0] main_bus_cti;
wire [1:0] main_bus_bte;
wire main_bus_err;
wire main_writer_sink_sink_stb;
reg main_writer_sink_sink_ack = 1'd1;
wire main_writer_sink_sink_eop;
wire [31:0] main_writer_sink_sink_payload_data;
wire [3:0] main_writer_sink_sink_payload_last_be;
wire [3:0] main_writer_sink_sink_payload_error;
wire [1:0] main_writer_slot_status;
wire [31:0] main_writer_length_status;
reg [31:0] main_writer_errors_status = 32'd0;
wire main_writer_irq;
wire main_writer_available_status;
wire main_writer_available_pending;
wire main_writer_available_trigger;
reg main_writer_available_clear;
wire main_writer_status_re;
wire main_writer_status_r;
wire main_writer_status_w;
wire main_writer_pending_re;
wire main_writer_pending_r;
wire main_writer_pending_w;
reg main_writer_storage_full = 1'd0;
wire main_writer_storage;
reg main_writer_re = 1'd0;
reg [2:0] main_writer_increment;
reg [31:0] main_writer_counter = 32'd0;
reg main_writer_counter_reset;
reg main_writer_counter_ce;
reg [1:0] main_writer_slot = 2'd0;
reg main_writer_slot_ce;
reg main_writer_ongoing;
reg main_writer_fifo_sink_stb;
wire main_writer_fifo_sink_ack;
reg main_writer_fifo_sink_eop = 1'd0;
wire [1:0] main_writer_fifo_sink_payload_slot;
wire [31:0] main_writer_fifo_sink_payload_length;
wire main_writer_fifo_source_stb;
wire main_writer_fifo_source_ack;
wire main_writer_fifo_source_eop;
wire [1:0] main_writer_fifo_source_payload_slot;
wire [31:0] main_writer_fifo_source_payload_length;
wire main_writer_fifo_syncfifo_we;
wire main_writer_fifo_syncfifo_writable;
wire main_writer_fifo_syncfifo_re;
wire main_writer_fifo_syncfifo_readable;
wire [34:0] main_writer_fifo_syncfifo_din;
wire [34:0] main_writer_fifo_syncfifo_dout;
reg [2:0] main_writer_fifo_level = 3'd0;
reg main_writer_fifo_replace = 1'd0;
reg [1:0] main_writer_fifo_produce = 2'd0;
reg [1:0] main_writer_fifo_consume = 2'd0;
reg [1:0] main_writer_fifo_wrport_adr;
wire [34:0] main_writer_fifo_wrport_dat_r;
wire main_writer_fifo_wrport_we;
wire [34:0] main_writer_fifo_wrport_dat_w;
wire main_writer_fifo_do_read;
wire [1:0] main_writer_fifo_rdport_adr;
wire [34:0] main_writer_fifo_rdport_dat_r;
wire [1:0] main_writer_fifo_fifo_in_payload_slot;
wire [31:0] main_writer_fifo_fifo_in_payload_length;
wire main_writer_fifo_fifo_in_eop;
wire [1:0] main_writer_fifo_fifo_out_payload_slot;
wire [31:0] main_writer_fifo_fifo_out_payload_length;
wire main_writer_fifo_fifo_out_eop;
reg [8:0] main_writer_memory0_adr;
wire [31:0] main_writer_memory0_dat_r;
reg main_writer_memory0_we;
reg [31:0] main_writer_memory0_dat_w;
reg [8:0] main_writer_memory1_adr;
wire [31:0] main_writer_memory1_dat_r;
reg main_writer_memory1_we;
reg [31:0] main_writer_memory1_dat_w;
reg [8:0] main_writer_memory2_adr;
wire [31:0] main_writer_memory2_dat_r;
reg main_writer_memory2_we;
reg [31:0] main_writer_memory2_dat_w;
reg [8:0] main_writer_memory3_adr;
wire [31:0] main_writer_memory3_dat_r;
reg main_writer_memory3_we;
reg [31:0] main_writer_memory3_dat_w;
reg main_reader_source_source_stb;
wire main_reader_source_source_ack;
reg main_reader_source_source_eop;
reg [31:0] main_reader_source_source_payload_data;
reg [3:0] main_reader_source_source_payload_last_be;
reg [3:0] main_reader_source_source_payload_error = 4'd0;
wire main_reader_start_re;
wire main_reader_start_r;
reg main_reader_start_w = 1'd0;
wire main_reader_ready_status;
reg [1:0] main_reader_slot_storage_full = 2'd0;
wire [1:0] main_reader_slot_storage;
reg main_reader_slot_re = 1'd0;
reg [10:0] main_reader_length_storage_full = 11'd0;
wire [10:0] main_reader_length_storage;
reg main_reader_length_re = 1'd0;
wire main_reader_irq;
wire main_reader_done_status;
reg main_reader_done_pending = 1'd0;
reg main_reader_done_trigger;
reg main_reader_done_clear;
wire main_reader_eventmanager_status_re;
wire main_reader_eventmanager_status_r;
wire main_reader_eventmanager_status_w;
wire main_reader_eventmanager_pending_re;
wire main_reader_eventmanager_pending_r;
wire main_reader_eventmanager_pending_w;
reg main_reader_eventmanager_storage_full = 1'd0;
wire main_reader_eventmanager_storage;
reg main_reader_eventmanager_re = 1'd0;
wire main_reader_fifo_sink_stb;
wire main_reader_fifo_sink_ack;
reg main_reader_fifo_sink_eop = 1'd0;
wire [1:0] main_reader_fifo_sink_payload_slot;
wire [10:0] main_reader_fifo_sink_payload_length;
wire main_reader_fifo_source_stb;
reg main_reader_fifo_source_ack;
wire main_reader_fifo_source_eop;
wire [1:0] main_reader_fifo_source_payload_slot;
wire [10:0] main_reader_fifo_source_payload_length;
wire main_reader_fifo_syncfifo_we;
wire main_reader_fifo_syncfifo_writable;
wire main_reader_fifo_syncfifo_re;
wire main_reader_fifo_syncfifo_readable;
wire [13:0] main_reader_fifo_syncfifo_din;
wire [13:0] main_reader_fifo_syncfifo_dout;
reg [2:0] main_reader_fifo_level = 3'd0;
reg main_reader_fifo_replace = 1'd0;
reg [1:0] main_reader_fifo_produce = 2'd0;
reg [1:0] main_reader_fifo_consume = 2'd0;
reg [1:0] main_reader_fifo_wrport_adr;
wire [13:0] main_reader_fifo_wrport_dat_r;
wire main_reader_fifo_wrport_we;
wire [13:0] main_reader_fifo_wrport_dat_w;
wire main_reader_fifo_do_read;
wire [1:0] main_reader_fifo_rdport_adr;
wire [13:0] main_reader_fifo_rdport_dat_r;
wire [1:0] main_reader_fifo_fifo_in_payload_slot;
wire [10:0] main_reader_fifo_fifo_in_payload_length;
wire main_reader_fifo_fifo_in_eop;
wire [1:0] main_reader_fifo_fifo_out_payload_slot;
wire [10:0] main_reader_fifo_fifo_out_payload_length;
wire main_reader_fifo_fifo_out_eop;
reg [10:0] main_reader_counter = 11'd0;
reg main_reader_counter_reset;
reg main_reader_counter_ce;
wire main_reader_last;
reg main_reader_last_d = 1'd0;
wire [8:0] main_reader_memory0_adr;
wire [31:0] main_reader_memory0_dat_r;
wire [8:0] main_reader_memory1_adr;
wire [31:0] main_reader_memory1_dat_r;
wire [8:0] main_reader_memory2_adr;
wire [31:0] main_reader_memory2_dat_r;
wire [8:0] main_reader_memory3_adr;
wire [31:0] main_reader_memory3_dat_r;
wire main_ev_irq;
wire [29:0] main_sram0_bus_adr0;
wire [31:0] main_sram0_bus_dat_w0;
wire [31:0] main_sram0_bus_dat_r0;
wire [3:0] main_sram0_bus_sel0;
wire main_sram0_bus_cyc0;
wire main_sram0_bus_stb0;
reg main_sram0_bus_ack0 = 1'd0;
wire main_sram0_bus_we0;
wire [2:0] main_sram0_bus_cti0;
wire [1:0] main_sram0_bus_bte0;
reg main_sram0_bus_err0 = 1'd0;
wire [8:0] main_sram0_adr0;
wire [31:0] main_sram0_dat_r0;
wire [29:0] main_sram1_bus_adr0;
wire [31:0] main_sram1_bus_dat_w0;
wire [31:0] main_sram1_bus_dat_r0;
wire [3:0] main_sram1_bus_sel0;
wire main_sram1_bus_cyc0;
wire main_sram1_bus_stb0;
reg main_sram1_bus_ack0 = 1'd0;
wire main_sram1_bus_we0;
wire [2:0] main_sram1_bus_cti0;
wire [1:0] main_sram1_bus_bte0;
reg main_sram1_bus_err0 = 1'd0;
wire [8:0] main_sram1_adr0;
wire [31:0] main_sram1_dat_r0;
wire [29:0] main_sram2_bus_adr0;
wire [31:0] main_sram2_bus_dat_w0;
wire [31:0] main_sram2_bus_dat_r0;
wire [3:0] main_sram2_bus_sel0;
wire main_sram2_bus_cyc0;
wire main_sram2_bus_stb0;
reg main_sram2_bus_ack0 = 1'd0;
wire main_sram2_bus_we0;
wire [2:0] main_sram2_bus_cti0;
wire [1:0] main_sram2_bus_bte0;
reg main_sram2_bus_err0 = 1'd0;
wire [8:0] main_sram2_adr0;
wire [31:0] main_sram2_dat_r0;
wire [29:0] main_sram3_bus_adr0;
wire [31:0] main_sram3_bus_dat_w0;
wire [31:0] main_sram3_bus_dat_r0;
wire [3:0] main_sram3_bus_sel0;
wire main_sram3_bus_cyc0;
wire main_sram3_bus_stb0;
reg main_sram3_bus_ack0 = 1'd0;
wire main_sram3_bus_we0;
wire [2:0] main_sram3_bus_cti0;
wire [1:0] main_sram3_bus_bte0;
reg main_sram3_bus_err0 = 1'd0;
wire [8:0] main_sram3_adr0;
wire [31:0] main_sram3_dat_r0;
wire [29:0] main_sram0_bus_adr1;
wire [31:0] main_sram0_bus_dat_w1;
wire [31:0] main_sram0_bus_dat_r1;
wire [3:0] main_sram0_bus_sel1;
wire main_sram0_bus_cyc1;
wire main_sram0_bus_stb1;
reg main_sram0_bus_ack1 = 1'd0;
wire main_sram0_bus_we1;
wire [2:0] main_sram0_bus_cti1;
wire [1:0] main_sram0_bus_bte1;
reg main_sram0_bus_err1 = 1'd0;
wire [8:0] main_sram0_adr1;
wire [31:0] main_sram0_dat_r1;
reg [3:0] main_sram0_we;
wire [31:0] main_sram0_dat_w;
wire [29:0] main_sram1_bus_adr1;
wire [31:0] main_sram1_bus_dat_w1;
wire [31:0] main_sram1_bus_dat_r1;
wire [3:0] main_sram1_bus_sel1;
wire main_sram1_bus_cyc1;
wire main_sram1_bus_stb1;
reg main_sram1_bus_ack1 = 1'd0;
wire main_sram1_bus_we1;
wire [2:0] main_sram1_bus_cti1;
wire [1:0] main_sram1_bus_bte1;
reg main_sram1_bus_err1 = 1'd0;
wire [8:0] main_sram1_adr1;
wire [31:0] main_sram1_dat_r1;
reg [3:0] main_sram1_we;
wire [31:0] main_sram1_dat_w;
wire [29:0] main_sram2_bus_adr1;
wire [31:0] main_sram2_bus_dat_w1;
wire [31:0] main_sram2_bus_dat_r1;
wire [3:0] main_sram2_bus_sel1;
wire main_sram2_bus_cyc1;
wire main_sram2_bus_stb1;
reg main_sram2_bus_ack1 = 1'd0;
wire main_sram2_bus_we1;
wire [2:0] main_sram2_bus_cti1;
wire [1:0] main_sram2_bus_bte1;
reg main_sram2_bus_err1 = 1'd0;
wire [8:0] main_sram2_adr1;
wire [31:0] main_sram2_dat_r1;
reg [3:0] main_sram2_we;
wire [31:0] main_sram2_dat_w;
wire [29:0] main_sram3_bus_adr1;
wire [31:0] main_sram3_bus_dat_w1;
wire [31:0] main_sram3_bus_dat_r1;
wire [3:0] main_sram3_bus_sel1;
wire main_sram3_bus_cyc1;
wire main_sram3_bus_stb1;
reg main_sram3_bus_ack1 = 1'd0;
wire main_sram3_bus_we1;
wire [2:0] main_sram3_bus_cti1;
wire [1:0] main_sram3_bus_bte1;
reg main_sram3_bus_err1 = 1'd0;
wire [8:0] main_sram3_adr1;
wire [31:0] main_sram3_dat_r1;
reg [3:0] main_sram3_we;
wire [31:0] main_sram3_dat_w;
reg [7:0] main_slave_sel;
reg [7:0] main_slave_sel_r = 8'd0;
reg main_kernel_cpu_storage_full = 1'd1;
wire main_kernel_cpu_storage;
reg main_kernel_cpu_re = 1'd0;
wire sys_kernel_clk;
wire sys_kernel_rst;
wire [29:0] main_kernel_cpu_ibus_adr;
wire [31:0] main_kernel_cpu_ibus_dat_w;
wire [31:0] main_kernel_cpu_ibus_dat_r;
wire [3:0] main_kernel_cpu_ibus_sel;
wire main_kernel_cpu_ibus_cyc;
wire main_kernel_cpu_ibus_stb;
wire main_kernel_cpu_ibus_ack;
wire main_kernel_cpu_ibus_we;
wire [2:0] main_kernel_cpu_ibus_cti;
wire [1:0] main_kernel_cpu_ibus_bte;
wire main_kernel_cpu_ibus_err;
wire [29:0] main_kernel_cpu_dbus_adr;
wire [31:0] main_kernel_cpu_dbus_dat_w;
wire [31:0] main_kernel_cpu_dbus_dat_r;
wire [3:0] main_kernel_cpu_dbus_sel;
wire main_kernel_cpu_dbus_cyc;
wire main_kernel_cpu_dbus_stb;
wire main_kernel_cpu_dbus_ack;
wire main_kernel_cpu_dbus_we;
wire [2:0] main_kernel_cpu_dbus_cti;
wire [1:0] main_kernel_cpu_dbus_bte;
wire main_kernel_cpu_dbus_err;
reg [31:0] main_kernel_cpu_interrupt = 32'd0;
wire [31:0] main_kernel_cpu_i_adr_o;
wire [31:0] main_kernel_cpu_d_adr_o;
wire [29:0] main_kernel_cpu_wb_sdram_adr;
wire [31:0] main_kernel_cpu_wb_sdram_dat_w;
wire [31:0] main_kernel_cpu_wb_sdram_dat_r;
wire [3:0] main_kernel_cpu_wb_sdram_sel;
wire main_kernel_cpu_wb_sdram_cyc;
wire main_kernel_cpu_wb_sdram_stb;
wire main_kernel_cpu_wb_sdram_ack;
wire main_kernel_cpu_wb_sdram_we;
wire [2:0] main_kernel_cpu_wb_sdram_cti;
wire [1:0] main_kernel_cpu_wb_sdram_bte;
wire main_kernel_cpu_wb_sdram_err;
wire [29:0] main_mailbox_i1_adr;
wire [31:0] main_mailbox_i1_dat_w;
reg [31:0] main_mailbox_i1_dat_r = 32'd0;
wire [3:0] main_mailbox_i1_sel;
wire main_mailbox_i1_cyc;
wire main_mailbox_i1_stb;
reg main_mailbox_i1_ack = 1'd0;
wire main_mailbox_i1_we;
wire [2:0] main_mailbox_i1_cti;
wire [1:0] main_mailbox_i1_bte;
reg main_mailbox_i1_err = 1'd0;
wire [29:0] main_mailbox_i2_adr;
wire [31:0] main_mailbox_i2_dat_w;
reg [31:0] main_mailbox_i2_dat_r = 32'd0;
wire [3:0] main_mailbox_i2_sel;
wire main_mailbox_i2_cyc;
wire main_mailbox_i2_stb;
reg main_mailbox_i2_ack = 1'd0;
wire main_mailbox_i2_we;
wire [2:0] main_mailbox_i2_cti;
wire [1:0] main_mailbox_i2_bte;
reg main_mailbox_i2_err = 1'd0;
reg [31:0] main_mailbox0 = 32'd0;
reg [31:0] main_mailbox1 = 32'd0;
reg [31:0] main_mailbox2 = 32'd0;
reg [7:0] main_add_identifier_storage_full = 8'd0;
wire [7:0] main_add_identifier_storage;
reg main_add_identifier_re = 1'd0;
wire [7:0] main_add_identifier_status;
wire [4:0] main_add_identifier_adr;
wire [7:0] main_add_identifier_dat_r;
reg [63:0] main_load_storage_full = 64'd0;
wire [63:0] main_load_storage;
reg main_load_re = 1'd0;
reg [63:0] main_reload_storage_full = 64'd0;
wire [63:0] main_reload_storage;
reg main_reload_re = 1'd0;
reg main_en_storage_full = 1'd0;
wire main_en_storage;
reg main_en_re = 1'd0;
wire main_update_value_re;
wire main_update_value_r;
reg main_update_value_w = 1'd0;
reg [63:0] main_value_status = 64'd0;
wire main_irq;
wire main_zero_status;
reg main_zero_pending = 1'd0;
wire main_zero_trigger;
reg main_zero_clear;
reg main_zero_old_trigger = 1'd0;
wire main_eventmanager_status_re;
wire main_eventmanager_status_r;
wire main_eventmanager_status_w;
wire main_eventmanager_pending_re;
wire main_eventmanager_pending_r;
wire main_eventmanager_pending_w;
reg main_eventmanager_storage_full = 1'd0;
wire main_eventmanager_storage;
reg main_eventmanager_re = 1'd0;
reg [63:0] main_value = 64'd0;
reg [1:0] main_leds_storage_full = 2'd0;
wire [1:0] main_leds_storage;
reg main_leds_re = 1'd0;
reg [1:0] main_i2c_status0;
reg [1:0] main_i2c_out_storage_full = 2'd0;
wire [1:0] main_i2c_out_storage;
reg main_i2c_out_re = 1'd0;
reg [1:0] main_i2c_oe_storage_full = 2'd0;
wire [1:0] main_i2c_oe_storage;
reg main_i2c_oe_re = 1'd0;
wire main_i2c_tstriple0_o;
wire main_i2c_tstriple0_oe;
wire main_i2c_tstriple0_i;
wire main_i2c_status1;
wire main_i2c_tstriple1_o;
wire main_i2c_tstriple1_oe;
wire main_i2c_tstriple1_i;
wire main_i2c_status2;
reg [7:0] main_output_8x0_o = 8'd0;
reg main_output_8x0_t_in = 1'd0;
wire main_output_8x0_t_out;
wire main_output_8x0_pad_o;
reg main_output_8x0_stb = 1'd0;
reg main_output_8x0_busy = 1'd0;
reg main_output_8x0_data = 1'd0;
reg [2:0] main_output_8x0_fine_ts = 3'd0;
wire main_output_8x0_override_en;
wire main_output_8x0_override_o;
reg main_output_8x0_previous_data = 1'd0;
reg [7:0] main_output_8x1_o = 8'd0;
reg main_output_8x1_t_in = 1'd0;
wire main_output_8x1_t_out;
wire main_output_8x1_pad_o;
reg main_output_8x1_stb = 1'd0;
reg main_output_8x1_busy = 1'd0;
reg main_output_8x1_data = 1'd0;
reg [2:0] main_output_8x1_fine_ts = 3'd0;
wire main_output_8x1_override_en;
wire main_output_8x1_override_o;
reg main_output_8x1_previous_data = 1'd0;
reg [7:0] main_output_8x2_o = 8'd0;
reg main_output_8x2_t_in = 1'd0;
wire main_output_8x2_t_out;
wire main_output_8x2_pad_o;
reg main_output_8x2_stb = 1'd0;
reg main_output_8x2_busy = 1'd0;
reg main_output_8x2_data = 1'd0;
reg [2:0] main_output_8x2_fine_ts = 3'd0;
wire main_output_8x2_override_en;
wire main_output_8x2_override_o;
reg main_output_8x2_previous_data = 1'd0;
reg [7:0] main_inout_8x0_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x0_serdes_i0;
wire main_inout_8x0_serdes_oe;
wire main_inout_8x0_serdes_pad_i0;
wire main_inout_8x0_serdes_pad_o0;
wire [7:0] main_inout_8x0_serdes_i1;
wire main_inout_8x0_serdes_pad_i1;
wire [7:0] main_inout_8x0_serdes_o1;
wire main_inout_8x0_serdes_t_in;
wire main_inout_8x0_serdes_t_out;
wire main_inout_8x0_serdes_pad_o1;
reg main_inout_8x0_inout_8x0_ointerface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_ointerface0_busy = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_data = 2'd0;
reg [1:0] main_inout_8x0_inout_8x0_ointerface0_address = 2'd0;
reg [2:0] main_inout_8x0_inout_8x0_ointerface0_fine_ts = 3'd0;
reg main_inout_8x0_inout_8x0_iinterface0_stb = 1'd0;
reg main_inout_8x0_inout_8x0_iinterface0_data = 1'd0;
reg [2:0] main_inout_8x0_inout_8x0_iinterface0_fine_ts = 3'd0;
wire main_inout_8x0_inout_8x0_override_en;
wire main_inout_8x0_inout_8x0_override_o;
wire main_inout_8x0_inout_8x0_override_oe;
(* dont_touch = "true" *) reg main_inout_8x0_inout_8x0_oe = 1'd0;
wire main_inout_8x0_inout_8x0_input_state;
reg main_inout_8x0_inout_8x0_previous_data = 1'd0;
reg main_inout_8x0_inout_8x0_oe_k = 1'd0;
reg [1:0] main_inout_8x0_inout_8x0_sensitivity = 2'd0;
reg main_inout_8x0_inout_8x0_sample = 1'd0;
reg main_inout_8x0_inout_8x0_i_d = 1'd0;
wire [7:0] main_inout_8x0_inout_8x0_i;
reg [2:0] main_inout_8x0_inout_8x0_o;
wire main_inout_8x0_inout_8x0_n;
reg [7:0] main_output_8x3_o = 8'd0;
reg main_output_8x3_t_in = 1'd0;
wire main_output_8x3_t_out;
wire main_output_8x3_pad_o;
reg main_output_8x3_stb = 1'd0;
reg main_output_8x3_busy = 1'd0;
reg main_output_8x3_data = 1'd0;
reg [2:0] main_output_8x3_fine_ts = 3'd0;
wire main_output_8x3_override_en;
wire main_output_8x3_override_o;
reg main_output_8x3_previous_data = 1'd0;
reg [7:0] main_output_8x4_o = 8'd0;
reg main_output_8x4_t_in = 1'd0;
wire main_output_8x4_t_out;
wire main_output_8x4_pad_o;
reg main_output_8x4_stb = 1'd0;
reg main_output_8x4_busy = 1'd0;
reg main_output_8x4_data = 1'd0;
reg [2:0] main_output_8x4_fine_ts = 3'd0;
wire main_output_8x4_override_en;
wire main_output_8x4_override_o;
reg main_output_8x4_previous_data = 1'd0;
reg [7:0] main_output_8x5_o = 8'd0;
reg main_output_8x5_t_in = 1'd0;
wire main_output_8x5_t_out;
wire main_output_8x5_pad_o;
reg main_output_8x5_stb = 1'd0;
reg main_output_8x5_busy = 1'd0;
reg main_output_8x5_data = 1'd0;
reg [2:0] main_output_8x5_fine_ts = 3'd0;
wire main_output_8x5_override_en;
wire main_output_8x5_override_o;
reg main_output_8x5_previous_data = 1'd0;
reg [7:0] main_inout_8x1_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x1_serdes_i0;
wire main_inout_8x1_serdes_oe;
wire main_inout_8x1_serdes_pad_i0;
wire main_inout_8x1_serdes_pad_o0;
wire [7:0] main_inout_8x1_serdes_i1;
wire main_inout_8x1_serdes_pad_i1;
wire [7:0] main_inout_8x1_serdes_o1;
wire main_inout_8x1_serdes_t_in;
wire main_inout_8x1_serdes_t_out;
wire main_inout_8x1_serdes_pad_o1;
reg main_inout_8x1_inout_8x1_ointerface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_ointerface1_busy = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_data = 2'd0;
reg [1:0] main_inout_8x1_inout_8x1_ointerface1_address = 2'd0;
reg [2:0] main_inout_8x1_inout_8x1_ointerface1_fine_ts = 3'd0;
reg main_inout_8x1_inout_8x1_iinterface1_stb = 1'd0;
reg main_inout_8x1_inout_8x1_iinterface1_data = 1'd0;
reg [2:0] main_inout_8x1_inout_8x1_iinterface1_fine_ts = 3'd0;
wire main_inout_8x1_inout_8x1_override_en;
wire main_inout_8x1_inout_8x1_override_o;
wire main_inout_8x1_inout_8x1_override_oe;
(* dont_touch = "true" *) reg main_inout_8x1_inout_8x1_oe = 1'd0;
wire main_inout_8x1_inout_8x1_input_state;
reg main_inout_8x1_inout_8x1_previous_data = 1'd0;
reg main_inout_8x1_inout_8x1_oe_k = 1'd0;
reg [1:0] main_inout_8x1_inout_8x1_sensitivity = 2'd0;
reg main_inout_8x1_inout_8x1_sample = 1'd0;
reg main_inout_8x1_inout_8x1_i_d = 1'd0;
wire [7:0] main_inout_8x1_inout_8x1_i;
reg [2:0] main_inout_8x1_inout_8x1_o;
wire main_inout_8x1_inout_8x1_n;
reg [7:0] main_output_8x6_o = 8'd0;
reg main_output_8x6_t_in = 1'd0;
wire main_output_8x6_t_out;
wire main_output_8x6_pad_o;
reg main_output_8x6_stb = 1'd0;
reg main_output_8x6_busy = 1'd0;
reg main_output_8x6_data = 1'd0;
reg [2:0] main_output_8x6_fine_ts = 3'd0;
wire main_output_8x6_override_en;
wire main_output_8x6_override_o;
reg main_output_8x6_previous_data = 1'd0;
reg [7:0] main_output_8x7_o = 8'd0;
reg main_output_8x7_t_in = 1'd0;
wire main_output_8x7_t_out;
wire main_output_8x7_pad_o;
reg main_output_8x7_stb = 1'd0;
reg main_output_8x7_busy = 1'd0;
reg main_output_8x7_data = 1'd0;
reg [2:0] main_output_8x7_fine_ts = 3'd0;
wire main_output_8x7_override_en;
wire main_output_8x7_override_o;
reg main_output_8x7_previous_data = 1'd0;
reg [7:0] main_output_8x8_o = 8'd0;
reg main_output_8x8_t_in = 1'd0;
wire main_output_8x8_t_out;
wire main_output_8x8_pad_o;
reg main_output_8x8_stb = 1'd0;
reg main_output_8x8_busy = 1'd0;
reg main_output_8x8_data = 1'd0;
reg [2:0] main_output_8x8_fine_ts = 3'd0;
wire main_output_8x8_override_en;
wire main_output_8x8_override_o;
reg main_output_8x8_previous_data = 1'd0;
reg [7:0] main_inout_8x2_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x2_serdes_i0;
wire main_inout_8x2_serdes_oe;
wire main_inout_8x2_serdes_pad_i0;
wire main_inout_8x2_serdes_pad_o0;
wire [7:0] main_inout_8x2_serdes_i1;
wire main_inout_8x2_serdes_pad_i1;
wire [7:0] main_inout_8x2_serdes_o1;
wire main_inout_8x2_serdes_t_in;
wire main_inout_8x2_serdes_t_out;
wire main_inout_8x2_serdes_pad_o1;
reg main_inout_8x2_inout_8x2_ointerface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_ointerface2_busy = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_data = 2'd0;
reg [1:0] main_inout_8x2_inout_8x2_ointerface2_address = 2'd0;
reg [2:0] main_inout_8x2_inout_8x2_ointerface2_fine_ts = 3'd0;
reg main_inout_8x2_inout_8x2_iinterface2_stb = 1'd0;
reg main_inout_8x2_inout_8x2_iinterface2_data = 1'd0;
reg [2:0] main_inout_8x2_inout_8x2_iinterface2_fine_ts = 3'd0;
wire main_inout_8x2_inout_8x2_override_en;
wire main_inout_8x2_inout_8x2_override_o;
wire main_inout_8x2_inout_8x2_override_oe;
(* dont_touch = "true" *) reg main_inout_8x2_inout_8x2_oe = 1'd0;
wire main_inout_8x2_inout_8x2_input_state;
reg main_inout_8x2_inout_8x2_previous_data = 1'd0;
reg main_inout_8x2_inout_8x2_oe_k = 1'd0;
reg [1:0] main_inout_8x2_inout_8x2_sensitivity = 2'd0;
reg main_inout_8x2_inout_8x2_sample = 1'd0;
reg main_inout_8x2_inout_8x2_i_d = 1'd0;
wire [7:0] main_inout_8x2_inout_8x2_i;
reg [2:0] main_inout_8x2_inout_8x2_o;
wire main_inout_8x2_inout_8x2_n;
reg [7:0] main_output_8x9_o = 8'd0;
reg main_output_8x9_t_in = 1'd0;
wire main_output_8x9_t_out;
wire main_output_8x9_pad_o;
reg main_output_8x9_stb = 1'd0;
reg main_output_8x9_busy = 1'd0;
reg main_output_8x9_data = 1'd0;
reg [2:0] main_output_8x9_fine_ts = 3'd0;
wire main_output_8x9_override_en;
wire main_output_8x9_override_o;
reg main_output_8x9_previous_data = 1'd0;
reg [7:0] main_output_8x10_o = 8'd0;
reg main_output_8x10_t_in = 1'd0;
wire main_output_8x10_t_out;
wire main_output_8x10_pad_o;
reg main_output_8x10_stb = 1'd0;
reg main_output_8x10_busy = 1'd0;
reg main_output_8x10_data = 1'd0;
reg [2:0] main_output_8x10_fine_ts = 3'd0;
wire main_output_8x10_override_en;
wire main_output_8x10_override_o;
reg main_output_8x10_previous_data = 1'd0;
reg [7:0] main_output_8x11_o = 8'd0;
reg main_output_8x11_t_in = 1'd0;
wire main_output_8x11_t_out;
wire main_output_8x11_pad_o;
reg main_output_8x11_stb = 1'd0;
reg main_output_8x11_busy = 1'd0;
reg main_output_8x11_data = 1'd0;
reg [2:0] main_output_8x11_fine_ts = 3'd0;
wire main_output_8x11_override_en;
wire main_output_8x11_override_o;
reg main_output_8x11_previous_data = 1'd0;
reg [7:0] main_inout_8x3_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x3_serdes_i0;
wire main_inout_8x3_serdes_oe;
wire main_inout_8x3_serdes_pad_i0;
wire main_inout_8x3_serdes_pad_o0;
wire [7:0] main_inout_8x3_serdes_i1;
wire main_inout_8x3_serdes_pad_i1;
wire [7:0] main_inout_8x3_serdes_o1;
wire main_inout_8x3_serdes_t_in;
wire main_inout_8x3_serdes_t_out;
wire main_inout_8x3_serdes_pad_o1;
reg main_inout_8x3_inout_8x3_ointerface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_ointerface3_busy = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_data = 2'd0;
reg [1:0] main_inout_8x3_inout_8x3_ointerface3_address = 2'd0;
reg [2:0] main_inout_8x3_inout_8x3_ointerface3_fine_ts = 3'd0;
reg main_inout_8x3_inout_8x3_iinterface3_stb = 1'd0;
reg main_inout_8x3_inout_8x3_iinterface3_data = 1'd0;
reg [2:0] main_inout_8x3_inout_8x3_iinterface3_fine_ts = 3'd0;
wire main_inout_8x3_inout_8x3_override_en;
wire main_inout_8x3_inout_8x3_override_o;
wire main_inout_8x3_inout_8x3_override_oe;
(* dont_touch = "true" *) reg main_inout_8x3_inout_8x3_oe = 1'd0;
wire main_inout_8x3_inout_8x3_input_state;
reg main_inout_8x3_inout_8x3_previous_data = 1'd0;
reg main_inout_8x3_inout_8x3_oe_k = 1'd0;
reg [1:0] main_inout_8x3_inout_8x3_sensitivity = 2'd0;
reg main_inout_8x3_inout_8x3_sample = 1'd0;
reg main_inout_8x3_inout_8x3_i_d = 1'd0;
wire [7:0] main_inout_8x3_inout_8x3_i;
reg [2:0] main_inout_8x3_inout_8x3_o;
wire main_inout_8x3_inout_8x3_n;
reg [7:0] main_inout_8x4_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x4_serdes_i0;
wire main_inout_8x4_serdes_oe;
wire main_inout_8x4_serdes_pad_i0;
wire main_inout_8x4_serdes_pad_o0;
wire [7:0] main_inout_8x4_serdes_i1;
wire main_inout_8x4_serdes_pad_i1;
wire [7:0] main_inout_8x4_serdes_o1;
wire main_inout_8x4_serdes_t_in;
wire main_inout_8x4_serdes_t_out;
wire main_inout_8x4_serdes_pad_o1;
reg main_inout_8x4_inout_8x4_ointerface4_stb = 1'd0;
reg main_inout_8x4_inout_8x4_ointerface4_busy = 1'd0;
reg [1:0] main_inout_8x4_inout_8x4_ointerface4_data = 2'd0;
reg [1:0] main_inout_8x4_inout_8x4_ointerface4_address = 2'd0;
reg [2:0] main_inout_8x4_inout_8x4_ointerface4_fine_ts = 3'd0;
reg main_inout_8x4_inout_8x4_iinterface4_stb = 1'd0;
reg main_inout_8x4_inout_8x4_iinterface4_data = 1'd0;
reg [2:0] main_inout_8x4_inout_8x4_iinterface4_fine_ts = 3'd0;
wire main_inout_8x4_inout_8x4_override_en;
wire main_inout_8x4_inout_8x4_override_o;
wire main_inout_8x4_inout_8x4_override_oe;
(* dont_touch = "true" *) reg main_inout_8x4_inout_8x4_oe = 1'd0;
wire main_inout_8x4_inout_8x4_input_state;
reg main_inout_8x4_inout_8x4_previous_data = 1'd0;
reg main_inout_8x4_inout_8x4_oe_k = 1'd0;
reg [1:0] main_inout_8x4_inout_8x4_sensitivity = 2'd0;
reg main_inout_8x4_inout_8x4_sample = 1'd0;
reg main_inout_8x4_inout_8x4_i_d = 1'd0;
wire [7:0] main_inout_8x4_inout_8x4_i;
reg [2:0] main_inout_8x4_inout_8x4_o;
wire main_inout_8x4_inout_8x4_n;
reg [7:0] main_inout_8x5_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x5_serdes_i0;
wire main_inout_8x5_serdes_oe;
wire main_inout_8x5_serdes_pad_i0;
wire main_inout_8x5_serdes_pad_o0;
wire [7:0] main_inout_8x5_serdes_i1;
wire main_inout_8x5_serdes_pad_i1;
wire [7:0] main_inout_8x5_serdes_o1;
wire main_inout_8x5_serdes_t_in;
wire main_inout_8x5_serdes_t_out;
wire main_inout_8x5_serdes_pad_o1;
reg main_inout_8x5_inout_8x5_ointerface5_stb = 1'd0;
reg main_inout_8x5_inout_8x5_ointerface5_busy = 1'd0;
reg [1:0] main_inout_8x5_inout_8x5_ointerface5_data = 2'd0;
reg [1:0] main_inout_8x5_inout_8x5_ointerface5_address = 2'd0;
reg [2:0] main_inout_8x5_inout_8x5_ointerface5_fine_ts = 3'd0;
reg main_inout_8x5_inout_8x5_iinterface5_stb = 1'd0;
reg main_inout_8x5_inout_8x5_iinterface5_data = 1'd0;
reg [2:0] main_inout_8x5_inout_8x5_iinterface5_fine_ts = 3'd0;
wire main_inout_8x5_inout_8x5_override_en;
wire main_inout_8x5_inout_8x5_override_o;
wire main_inout_8x5_inout_8x5_override_oe;
(* dont_touch = "true" *) reg main_inout_8x5_inout_8x5_oe = 1'd0;
wire main_inout_8x5_inout_8x5_input_state;
reg main_inout_8x5_inout_8x5_previous_data = 1'd0;
reg main_inout_8x5_inout_8x5_oe_k = 1'd0;
reg [1:0] main_inout_8x5_inout_8x5_sensitivity = 2'd0;
reg main_inout_8x5_inout_8x5_sample = 1'd0;
reg main_inout_8x5_inout_8x5_i_d = 1'd0;
wire [7:0] main_inout_8x5_inout_8x5_i;
reg [2:0] main_inout_8x5_inout_8x5_o;
wire main_inout_8x5_inout_8x5_n;
reg [7:0] main_inout_8x6_serdes_o0 = 8'd0;
wire [7:0] main_inout_8x6_serdes_i0;
wire main_inout_8x6_serdes_oe;
wire main_inout_8x6_serdes_pad_i0;
wire main_inout_8x6_serdes_pad_o0;
wire [7:0] main_inout_8x6_serdes_i1;
wire main_inout_8x6_serdes_pad_i1;
wire [7:0] main_inout_8x6_serdes_o1;
wire main_inout_8x6_serdes_t_in;
wire main_inout_8x6_serdes_t_out;
wire main_inout_8x6_serdes_pad_o1;
reg main_inout_8x6_inout_8x6_ointerface6_stb = 1'd0;
reg main_inout_8x6_inout_8x6_ointerface6_busy = 1'd0;
reg [1:0] main_inout_8x6_inout_8x6_ointerface6_data = 2'd0;
reg [1:0] main_inout_8x6_inout_8x6_ointerface6_address = 2'd0;
reg [2:0] main_inout_8x6_inout_8x6_ointerface6_fine_ts = 3'd0;
reg main_inout_8x6_inout_8x6_iinterface6_stb = 1'd0;
reg main_inout_8x6_inout_8x6_iinterface6_data = 1'd0;
reg [2:0] main_inout_8x6_inout_8x6_iinterface6_fine_ts = 3'd0;
wire main_inout_8x6_inout_8x6_override_en;
wire main_inout_8x6_inout_8x6_override_o;
wire main_inout_8x6_inout_8x6_override_oe;
(* dont_touch = "true" *) reg main_inout_8x6_inout_8x6_oe = 1'd0;
wire main_inout_8x6_inout_8x6_input_state;
reg main_inout_8x6_inout_8x6_previous_data = 1'd0;
reg main_inout_8x6_inout_8x6_oe_k = 1'd0;
reg [1:0] main_inout_8x6_inout_8x6_sensitivity = 2'd0;
reg main_inout_8x6_inout_8x6_sample = 1'd0;
reg main_inout_8x6_inout_8x6_i_d = 1'd0;
wire [7:0] main_inout_8x6_inout_8x6_i;
reg [2:0] main_inout_8x6_inout_8x6_o;
wire main_inout_8x6_inout_8x6_n;
reg main_output0_stb = 1'd0;
reg main_output0_busy = 1'd0;
reg main_output0_data = 1'd0;
reg main_output0_pad_o = 1'd0;
wire main_output0_override_en;
wire main_output0_override_o;
reg main_output0_pad_k = 1'd0;
reg main_output1_stb = 1'd0;
reg main_output1_busy = 1'd0;
reg main_output1_data = 1'd0;
reg main_output1_pad_o = 1'd0;
wire main_output1_override_en;
wire main_output1_override_o;
reg main_output1_pad_k = 1'd0;
reg main_clockgen_stb = 1'd0;
reg main_clockgen_busy = 1'd0;
reg [23:0] main_clockgen_data = 24'd0;
reg [23:0] main_clockgen_ftw = 24'd0;
reg [23:0] main_clockgen_acc = 24'd0;
wire main_spimaster0_interface_cs;
wire main_spimaster0_interface_cs_polarity;
wire main_spimaster0_interface_clk_next;
wire main_spimaster0_interface_clk_polarity;
wire main_spimaster0_interface_cs_next;
wire main_spimaster0_interface_ce;
wire main_spimaster0_interface_sample;
wire main_spimaster0_interface_offline;
wire main_spimaster0_interface_half_duplex;
reg main_spimaster0_interface_sdi;
wire main_spimaster0_interface_sdo;
reg main_spimaster0_interface_cs_o = 1'd1;
wire main_spimaster0_interface_cs_oe;
wire main_spimaster0_interface_cs_i;
reg main_spimaster0_interface_clk_o = 1'd0;
wire main_spimaster0_interface_clk_oe;
wire main_spimaster0_interface_clk_i;
wire main_spimaster0_interface_mosi_o;
wire main_spimaster0_interface_mosi_oe;
wire main_spimaster0_interface_mosi_i;
wire main_spimaster0_interface_miso_o;
wire main_spimaster0_interface_miso_oe;
reg main_spimaster0_interface_miso_i = 1'd0;
reg main_spimaster0_interface_miso_reg = 1'd0;
reg main_spimaster0_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster0_spimachine0_length;
wire main_spimaster0_spimachine0_clk_phase;
reg main_spimaster0_spimachine0_clk_next;
reg main_spimaster0_spimachine0_cs_next;
wire main_spimaster0_spimachine0_ce;
reg main_spimaster0_spimachine0_idle;
wire main_spimaster0_spimachine0_load0;
reg main_spimaster0_spimachine0_readable;
reg main_spimaster0_spimachine0_writable;
wire main_spimaster0_spimachine0_end0;
wire [31:0] main_spimaster0_spimachine0_pdo;
wire [31:0] main_spimaster0_spimachine0_pdi;
reg main_spimaster0_spimachine0_sdo = 1'd0;
wire main_spimaster0_spimachine0_sdi;
wire main_spimaster0_spimachine0_lsb_first;
reg main_spimaster0_spimachine0_load1;
reg main_spimaster0_spimachine0_shift;
reg main_spimaster0_spimachine0_sample;
reg [31:0] main_spimaster0_spimachine0_sr = 32'd0;
wire [7:0] main_spimaster0_spimachine0_div;
reg main_spimaster0_spimachine0_extend;
wire main_spimaster0_spimachine0_done;
reg main_spimaster0_spimachine0_count;
reg [6:0] main_spimaster0_spimachine0_cnt = 7'd0;
wire main_spimaster0_spimachine0_cnt_done;
reg main_spimaster0_spimachine0_do_extend = 1'd0;
reg [4:0] main_spimaster0_spimachine0_n = 5'd0;
reg main_spimaster0_spimachine0_end1 = 1'd0;
reg main_spimaster0_ointerface0_stb = 1'd0;
wire main_spimaster0_ointerface0_busy;
reg [31:0] main_spimaster0_ointerface0_data = 32'd0;
reg main_spimaster0_ointerface0_address = 1'd0;
wire main_spimaster0_iinterface0_stb;
wire [31:0] main_spimaster0_iinterface0_data;
reg main_spimaster0_config_offline = 1'd1;
reg main_spimaster0_config_end = 1'd1;
reg main_spimaster0_config_input = 1'd0;
reg main_spimaster0_config_cs_polarity = 1'd0;
reg main_spimaster0_config_clk_polarity = 1'd0;
reg main_spimaster0_config_clk_phase = 1'd0;
reg main_spimaster0_config_lsb_first = 1'd0;
reg main_spimaster0_config_half_duplex = 1'd0;
reg [4:0] main_spimaster0_config_length = 5'd0;
reg [2:0] main_spimaster0_config_padding = 3'd0;
reg [7:0] main_spimaster0_config_div = 8'd0;
reg [7:0] main_spimaster0_config_cs = 8'd0;
reg main_spimaster0_read = 1'd0;
wire main_spimaster1_interface_cs;
wire main_spimaster1_interface_cs_polarity;
wire main_spimaster1_interface_clk_next;
wire main_spimaster1_interface_clk_polarity;
wire main_spimaster1_interface_cs_next;
wire main_spimaster1_interface_ce;
wire main_spimaster1_interface_sample;
wire main_spimaster1_interface_offline;
wire main_spimaster1_interface_half_duplex;
reg main_spimaster1_interface_sdi;
wire main_spimaster1_interface_sdo;
reg main_spimaster1_interface_cs_o = 1'd1;
wire main_spimaster1_interface_cs_oe;
wire main_spimaster1_interface_cs_i;
reg main_spimaster1_interface_clk_o = 1'd0;
wire main_spimaster1_interface_clk_oe;
wire main_spimaster1_interface_clk_i;
wire main_spimaster1_interface_mosi_o;
wire main_spimaster1_interface_mosi_oe;
wire main_spimaster1_interface_mosi_i;
wire main_spimaster1_interface_miso_o;
wire main_spimaster1_interface_miso_oe;
wire main_spimaster1_interface_miso_i;
reg main_spimaster1_interface_miso_reg = 1'd0;
reg main_spimaster1_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster1_spimachine1_length;
wire main_spimaster1_spimachine1_clk_phase;
reg main_spimaster1_spimachine1_clk_next;
reg main_spimaster1_spimachine1_cs_next;
wire main_spimaster1_spimachine1_ce;
reg main_spimaster1_spimachine1_idle;
wire main_spimaster1_spimachine1_load0;
reg main_spimaster1_spimachine1_readable;
reg main_spimaster1_spimachine1_writable;
wire main_spimaster1_spimachine1_end0;
wire [31:0] main_spimaster1_spimachine1_pdo;
wire [31:0] main_spimaster1_spimachine1_pdi;
reg main_spimaster1_spimachine1_sdo = 1'd0;
wire main_spimaster1_spimachine1_sdi;
wire main_spimaster1_spimachine1_lsb_first;
reg main_spimaster1_spimachine1_load1;
reg main_spimaster1_spimachine1_shift;
reg main_spimaster1_spimachine1_sample;
reg [31:0] main_spimaster1_spimachine1_sr = 32'd0;
wire [7:0] main_spimaster1_spimachine1_div;
reg main_spimaster1_spimachine1_extend;
wire main_spimaster1_spimachine1_done;
reg main_spimaster1_spimachine1_count;
reg [6:0] main_spimaster1_spimachine1_cnt = 7'd0;
wire main_spimaster1_spimachine1_cnt_done;
reg main_spimaster1_spimachine1_do_extend = 1'd0;
reg [4:0] main_spimaster1_spimachine1_n = 5'd0;
reg main_spimaster1_spimachine1_end1 = 1'd0;
reg main_spimaster1_ointerface1_stb = 1'd0;
wire main_spimaster1_ointerface1_busy;
reg [31:0] main_spimaster1_ointerface1_data = 32'd0;
reg main_spimaster1_ointerface1_address = 1'd0;
wire main_spimaster1_iinterface1_stb;
wire [31:0] main_spimaster1_iinterface1_data;
reg main_spimaster1_config_offline = 1'd1;
reg main_spimaster1_config_end = 1'd1;
reg main_spimaster1_config_input = 1'd0;
reg main_spimaster1_config_cs_polarity = 1'd0;
reg main_spimaster1_config_clk_polarity = 1'd0;
reg main_spimaster1_config_clk_phase = 1'd0;
reg main_spimaster1_config_lsb_first = 1'd0;
reg main_spimaster1_config_half_duplex = 1'd0;
reg [4:0] main_spimaster1_config_length = 5'd0;
reg [2:0] main_spimaster1_config_padding = 3'd0;
reg [7:0] main_spimaster1_config_div = 8'd0;
reg [7:0] main_spimaster1_config_cs = 8'd0;
reg main_spimaster1_read = 1'd0;
wire main_spimaster2_interface_cs;
wire main_spimaster2_interface_cs_polarity;
wire main_spimaster2_interface_clk_next;
wire main_spimaster2_interface_clk_polarity;
wire main_spimaster2_interface_cs_next;
wire main_spimaster2_interface_ce;
wire main_spimaster2_interface_sample;
wire main_spimaster2_interface_offline;
wire main_spimaster2_interface_half_duplex;
reg main_spimaster2_interface_sdi;
wire main_spimaster2_interface_sdo;
reg main_spimaster2_interface_cs_o = 1'd1;
wire main_spimaster2_interface_cs_oe;
wire main_spimaster2_interface_cs_i;
reg main_spimaster2_interface_clk_o = 1'd0;
wire main_spimaster2_interface_clk_oe;
wire main_spimaster2_interface_clk_i;
wire main_spimaster2_interface_mosi_o;
wire main_spimaster2_interface_mosi_oe;
wire main_spimaster2_interface_mosi_i;
wire main_spimaster2_interface_miso_o;
wire main_spimaster2_interface_miso_oe;
wire main_spimaster2_interface_miso_i;
reg main_spimaster2_interface_miso_reg = 1'd0;
reg main_spimaster2_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster2_spimachine2_length;
wire main_spimaster2_spimachine2_clk_phase;
reg main_spimaster2_spimachine2_clk_next;
reg main_spimaster2_spimachine2_cs_next;
wire main_spimaster2_spimachine2_ce;
reg main_spimaster2_spimachine2_idle;
wire main_spimaster2_spimachine2_load0;
reg main_spimaster2_spimachine2_readable;
reg main_spimaster2_spimachine2_writable;
wire main_spimaster2_spimachine2_end0;
wire [31:0] main_spimaster2_spimachine2_pdo;
wire [31:0] main_spimaster2_spimachine2_pdi;
reg main_spimaster2_spimachine2_sdo = 1'd0;
wire main_spimaster2_spimachine2_sdi;
wire main_spimaster2_spimachine2_lsb_first;
reg main_spimaster2_spimachine2_load1;
reg main_spimaster2_spimachine2_shift;
reg main_spimaster2_spimachine2_sample;
reg [31:0] main_spimaster2_spimachine2_sr = 32'd0;
wire [7:0] main_spimaster2_spimachine2_div;
reg main_spimaster2_spimachine2_extend;
wire main_spimaster2_spimachine2_done;
reg main_spimaster2_spimachine2_count;
reg [6:0] main_spimaster2_spimachine2_cnt = 7'd0;
wire main_spimaster2_spimachine2_cnt_done;
reg main_spimaster2_spimachine2_do_extend = 1'd0;
reg [4:0] main_spimaster2_spimachine2_n = 5'd0;
reg main_spimaster2_spimachine2_end1 = 1'd0;
reg main_spimaster2_ointerface2_stb = 1'd0;
wire main_spimaster2_ointerface2_busy;
reg [31:0] main_spimaster2_ointerface2_data = 32'd0;
reg main_spimaster2_ointerface2_address = 1'd0;
wire main_spimaster2_iinterface2_stb;
wire [31:0] main_spimaster2_iinterface2_data;
reg main_spimaster2_config_offline = 1'd1;
reg main_spimaster2_config_end = 1'd1;
reg main_spimaster2_config_input = 1'd0;
reg main_spimaster2_config_cs_polarity = 1'd0;
reg main_spimaster2_config_clk_polarity = 1'd0;
reg main_spimaster2_config_clk_phase = 1'd0;
reg main_spimaster2_config_lsb_first = 1'd0;
reg main_spimaster2_config_half_duplex = 1'd0;
reg [4:0] main_spimaster2_config_length = 5'd0;
reg [2:0] main_spimaster2_config_padding = 3'd0;
reg [7:0] main_spimaster2_config_div = 8'd0;
reg [7:0] main_spimaster2_config_cs = 8'd0;
reg main_spimaster2_read = 1'd0;
wire main_spimaster3_interface_cs;
wire main_spimaster3_interface_cs_polarity;
wire main_spimaster3_interface_clk_next;
wire main_spimaster3_interface_clk_polarity;
wire main_spimaster3_interface_cs_next;
wire main_spimaster3_interface_ce;
wire main_spimaster3_interface_sample;
wire main_spimaster3_interface_offline;
wire main_spimaster3_interface_half_duplex;
reg main_spimaster3_interface_sdi;
wire main_spimaster3_interface_sdo;
reg main_spimaster3_interface_cs_o = 1'd1;
wire main_spimaster3_interface_cs_oe;
wire main_spimaster3_interface_cs_i;
reg main_spimaster3_interface_clk_o = 1'd0;
wire main_spimaster3_interface_clk_oe;
wire main_spimaster3_interface_clk_i;
wire main_spimaster3_interface_mosi_o;
wire main_spimaster3_interface_mosi_oe;
wire main_spimaster3_interface_mosi_i;
wire main_spimaster3_interface_miso_o;
wire main_spimaster3_interface_miso_oe;
wire main_spimaster3_interface_miso_i;
reg main_spimaster3_interface_miso_reg = 1'd0;
reg main_spimaster3_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster3_spimachine3_length;
wire main_spimaster3_spimachine3_clk_phase;
reg main_spimaster3_spimachine3_clk_next;
reg main_spimaster3_spimachine3_cs_next;
wire main_spimaster3_spimachine3_ce;
reg main_spimaster3_spimachine3_idle;
wire main_spimaster3_spimachine3_load0;
reg main_spimaster3_spimachine3_readable;
reg main_spimaster3_spimachine3_writable;
wire main_spimaster3_spimachine3_end0;
wire [31:0] main_spimaster3_spimachine3_pdo;
wire [31:0] main_spimaster3_spimachine3_pdi;
reg main_spimaster3_spimachine3_sdo = 1'd0;
wire main_spimaster3_spimachine3_sdi;
wire main_spimaster3_spimachine3_lsb_first;
reg main_spimaster3_spimachine3_load1;
reg main_spimaster3_spimachine3_shift;
reg main_spimaster3_spimachine3_sample;
reg [31:0] main_spimaster3_spimachine3_sr = 32'd0;
wire [7:0] main_spimaster3_spimachine3_div;
reg main_spimaster3_spimachine3_extend;
wire main_spimaster3_spimachine3_done;
reg main_spimaster3_spimachine3_count;
reg [6:0] main_spimaster3_spimachine3_cnt = 7'd0;
wire main_spimaster3_spimachine3_cnt_done;
reg main_spimaster3_spimachine3_do_extend = 1'd0;
reg [4:0] main_spimaster3_spimachine3_n = 5'd0;
reg main_spimaster3_spimachine3_end1 = 1'd0;
reg main_spimaster3_ointerface3_stb = 1'd0;
wire main_spimaster3_ointerface3_busy;
reg [31:0] main_spimaster3_ointerface3_data = 32'd0;
reg main_spimaster3_ointerface3_address = 1'd0;
wire main_spimaster3_iinterface3_stb;
wire [31:0] main_spimaster3_iinterface3_data;
reg main_spimaster3_config_offline = 1'd1;
reg main_spimaster3_config_end = 1'd1;
reg main_spimaster3_config_input = 1'd0;
reg main_spimaster3_config_cs_polarity = 1'd0;
reg main_spimaster3_config_clk_polarity = 1'd0;
reg main_spimaster3_config_clk_phase = 1'd0;
reg main_spimaster3_config_lsb_first = 1'd0;
reg main_spimaster3_config_half_duplex = 1'd0;
reg [4:0] main_spimaster3_config_length = 5'd0;
reg [2:0] main_spimaster3_config_padding = 3'd0;
reg [7:0] main_spimaster3_config_div = 8'd0;
reg [7:0] main_spimaster3_config_cs = 8'd0;
reg main_spimaster3_read = 1'd0;
wire main_spimaster4_interface_cs;
wire main_spimaster4_interface_cs_polarity;
wire main_spimaster4_interface_clk_next;
wire main_spimaster4_interface_clk_polarity;
wire main_spimaster4_interface_cs_next;
wire main_spimaster4_interface_ce;
wire main_spimaster4_interface_sample;
wire main_spimaster4_interface_offline;
wire main_spimaster4_interface_half_duplex;
reg main_spimaster4_interface_sdi;
wire main_spimaster4_interface_sdo;
reg main_spimaster4_interface_cs_o = 1'd1;
wire main_spimaster4_interface_cs_oe;
wire main_spimaster4_interface_cs_i;
reg main_spimaster4_interface_clk_o = 1'd0;
wire main_spimaster4_interface_clk_oe;
wire main_spimaster4_interface_clk_i;
wire main_spimaster4_interface_mosi_o;
wire main_spimaster4_interface_mosi_oe;
wire main_spimaster4_interface_mosi_i;
wire main_spimaster4_interface_miso_o;
wire main_spimaster4_interface_miso_oe;
wire main_spimaster4_interface_miso_i;
reg main_spimaster4_interface_miso_reg = 1'd0;
reg main_spimaster4_interface_mosi_reg = 1'd0;
wire [4:0] main_spimaster4_spimachine4_length;
wire main_spimaster4_spimachine4_clk_phase;
reg main_spimaster4_spimachine4_clk_next;
reg main_spimaster4_spimachine4_cs_next;
wire main_spimaster4_spimachine4_ce;
reg main_spimaster4_spimachine4_idle;
wire main_spimaster4_spimachine4_load0;
reg main_spimaster4_spimachine4_readable;
reg main_spimaster4_spimachine4_writable;
wire main_spimaster4_spimachine4_end0;
wire [31:0] main_spimaster4_spimachine4_pdo;
wire [31:0] main_spimaster4_spimachine4_pdi;
reg main_spimaster4_spimachine4_sdo = 1'd0;
wire main_spimaster4_spimachine4_sdi;
wire main_spimaster4_spimachine4_lsb_first;
reg main_spimaster4_spimachine4_load1;
reg main_spimaster4_spimachine4_shift;
reg main_spimaster4_spimachine4_sample;
reg [31:0] main_spimaster4_spimachine4_sr = 32'd0;
wire [7:0] main_spimaster4_spimachine4_div;
reg main_spimaster4_spimachine4_extend;
wire main_spimaster4_spimachine4_done;
reg main_spimaster4_spimachine4_count;
reg [6:0] main_spimaster4_spimachine4_cnt = 7'd0;
wire main_spimaster4_spimachine4_cnt_done;
reg main_spimaster4_spimachine4_do_extend = 1'd0;
reg [4:0] main_spimaster4_spimachine4_n = 5'd0;
reg main_spimaster4_spimachine4_end1 = 1'd0;
reg main_spimaster4_ointerface4_stb = 1'd0;
wire main_spimaster4_ointerface4_busy;
reg [31:0] main_spimaster4_ointerface4_data = 32'd0;
reg main_spimaster4_ointerface4_address = 1'd0;
wire main_spimaster4_iinterface4_stb;
wire [31:0] main_spimaster4_iinterface4_data;
reg main_spimaster4_config_offline = 1'd1;
reg main_spimaster4_config_end = 1'd1;
reg main_spimaster4_config_input = 1'd0;
reg main_spimaster4_config_cs_polarity = 1'd0;
reg main_spimaster4_config_clk_polarity = 1'd0;
reg main_spimaster4_config_clk_phase = 1'd0;
reg main_spimaster4_config_lsb_first = 1'd0;
reg main_spimaster4_config_half_duplex = 1'd0;
reg [4:0] main_spimaster4_config_length = 5'd0;
reg [2:0] main_spimaster4_config_padding = 3'd0;
reg [7:0] main_spimaster4_config_div = 8'd0;
reg [7:0] main_spimaster4_config_cs = 8'd0;
reg main_spimaster4_read = 1'd0;
reg [29:0] main_ad9914_bus_adr = 30'd0;
reg [15:0] main_ad9914_bus_dat_w = 16'd0;
reg [15:0] main_ad9914_bus_dat_r;
reg [1:0] main_ad9914_bus_sel = 2'd0;
wire main_ad9914_bus_cyc;
wire main_ad9914_bus_stb;
reg main_ad9914_bus_ack;
reg main_ad9914_bus_we = 1'd0;
reg [15:0] main_ad9914_o = 16'd0;
reg main_ad9914_oe = 1'd0;
wire [15:0] main_ad9914_i;
reg main_ad9914_hold_address;
reg [15:0] main_ad9914_dr = 16'd0;
reg main_ad9914_rx;
reg [11:0] main_ad9914_gpio = 12'd0;
reg main_ad9914_gpio_load;
reg main_ad9914_bus_r_gpio;
reg main_ad9914_fud;
reg main_ad9914_wr;
reg main_ad9914_rd;
reg main_ad9914_read_timer_wait;
wire main_ad9914_read_timer_done;
reg [3:0] main_ad9914_read_timer_count = 4'd10;
reg main_ad9914_hiz_timer_wait;
wire main_ad9914_hiz_timer_done;
reg [1:0] main_ad9914_hiz_timer_count = 2'd3;
reg main_ad9914_stb = 1'd0;
wire main_ad9914_busy;
reg [15:0] main_ad9914_data = 16'd0;
reg [7:0] main_ad9914_address = 8'd0;
reg main_ad9914_active = 1'd0;
reg [31:0] main_ad9914_probes0 = 32'd0;
reg [31:0] main_ad9914_probes1 = 32'd0;
reg [31:0] main_ad9914_probes2 = 32'd0;
reg [31:0] main_ad9914_probes3 = 32'd0;
reg [31:0] main_ad9914_probes4 = 32'd0;
reg [31:0] main_ad9914_probes5 = 32'd0;
reg [31:0] main_ad9914_probes6 = 32'd0;
reg [31:0] main_ad9914_probes7 = 32'd0;
reg [31:0] main_ad9914_probes8 = 32'd0;
reg [31:0] main_ad9914_probes9 = 32'd0;
reg [31:0] main_ad9914_probes10 = 32'd0;
reg [7:0] main_ad9914_current_address = 8'd0;
reg [15:0] main_ad9914_current_data = 16'd0;
reg [14:0] main_ad9914_current_sel = 15'd0;
reg [31:0] main_ad9914_ftws0 = 32'd0;
reg [31:0] main_ad9914_ftws1 = 32'd0;
reg [31:0] main_ad9914_ftws2 = 32'd0;
reg [31:0] main_ad9914_ftws3 = 32'd0;
reg [31:0] main_ad9914_ftws4 = 32'd0;
reg [31:0] main_ad9914_ftws5 = 32'd0;
reg [31:0] main_ad9914_ftws6 = 32'd0;
reg [31:0] main_ad9914_ftws7 = 32'd0;
reg [31:0] main_ad9914_ftws8 = 32'd0;
reg [31:0] main_ad9914_ftws9 = 32'd0;
reg [31:0] main_ad9914_ftws10 = 32'd0;
reg main_stb = 1'd0;
reg main_busy = 1'd0;
reg [31:0] main_data = 32'd0;
reg main_rtio_crg_clock_sel_storage_full = 1'd0;
wire main_rtio_crg_clock_sel_storage;
reg main_rtio_crg_clock_sel_re = 1'd0;
reg main_rtio_crg_pll_reset_storage_full = 1'd1;
wire main_rtio_crg_pll_reset_storage;
reg main_rtio_crg_pll_reset_re = 1'd0;
wire main_rtio_crg_pll_locked_status;
wire rtio_clk;
wire rtio_rst;
wire rtiox4_clk;
wire ext_clkout_clk;
wire main_rtio_crg_rtio_external_clk;
wire main_rtio_crg_pll_locked;
wire main_rtio_crg_rtio_clk;
wire main_rtio_crg_rtiox4_clk;
wire main_rtio_crg_ext_clkout_clk;
reg [60:0] main_coarse_ts = 61'd0;
wire [63:0] main_full_ts;
wire [60:0] main_coarse_ts_sys;
wire [63:0] main_full_ts_sys;
reg main_load = 1'd0;
reg [60:0] main_load_value = 61'd0;
wire [60:0] main_i;
reg [60:0] main_o = 61'd0;
(* dont_touch = "true" *) reg [60:0] main_value_gray_rtio = 61'd0;
wire [60:0] main_value_gray_sys;
reg [60:0] main_value_sys;
reg [1:0] main_rtio_core_cri_cmd;
wire [23:0] main_rtio_core_cri_chan_sel;
wire [63:0] main_rtio_core_cri_o_timestamp;
wire [511:0] main_rtio_core_cri_o_data;
wire [7:0] main_rtio_core_cri_o_address;
wire [2:0] main_rtio_core_cri_o_status;
reg main_rtio_core_cri_o_buffer_space_valid = 1'd0;
reg [15:0] main_rtio_core_cri_o_buffer_space = 16'd0;
wire [63:0] main_rtio_core_cri_i_timeout;
reg [31:0] main_rtio_core_cri_i_data = 32'd0;
reg [63:0] main_rtio_core_cri_i_timestamp = 64'd0;
reg [3:0] main_rtio_core_cri_i_status = 4'd0;
wire main_rtio_core_reset_re;
wire main_rtio_core_reset_r;
reg main_rtio_core_reset_w = 1'd0;
wire main_rtio_core_reset_phy_re;
wire main_rtio_core_reset_phy_r;
reg main_rtio_core_reset_phy_w = 1'd0;
wire main_rtio_core_async_error_re;
wire [2:0] main_rtio_core_async_error_r;
wire [2:0] main_rtio_core_async_error_w;
reg [15:0] main_rtio_core_collision_channel_status = 16'd0;
reg [15:0] main_rtio_core_busy_channel_status = 16'd0;
reg [15:0] main_rtio_core_sequence_error_channel_status = 16'd0;
(* dont_touch = "true" *) reg main_rtio_core_cmd_reset = 1'd1;
(* dont_touch = "true" *) reg main_rtio_core_cmd_reset_phy = 1'd1;
wire rsys_clk;
wire rsys_rst;
wire rio_clk;
wire rio_rst;
wire rio_phy_clk;
wire rio_phy_rst;
reg main_rtio_core_outputs_lanedistributor_sequence_error = 1'd0;
reg [15:0] main_rtio_core_outputs_lanedistributor_sequence_error_channel = 16'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp = 61'd0;
reg main_rtio_core_outputs_lanedistributor_record0_we;
wire main_rtio_core_outputs_lanedistributor_record0_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record0_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record0_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record0_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record0_payload_data;
reg main_rtio_core_outputs_lanedistributor_record1_we;
wire main_rtio_core_outputs_lanedistributor_record1_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record1_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record1_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record1_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record1_payload_data;
reg main_rtio_core_outputs_lanedistributor_record2_we;
wire main_rtio_core_outputs_lanedistributor_record2_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record2_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record2_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record2_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record2_payload_data;
reg main_rtio_core_outputs_lanedistributor_record3_we;
wire main_rtio_core_outputs_lanedistributor_record3_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record3_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record3_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record3_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record3_payload_data;
reg main_rtio_core_outputs_lanedistributor_record4_we;
wire main_rtio_core_outputs_lanedistributor_record4_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record4_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record4_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record4_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record4_payload_data;
reg main_rtio_core_outputs_lanedistributor_record5_we;
wire main_rtio_core_outputs_lanedistributor_record5_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record5_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record5_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record5_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record5_payload_data;
reg main_rtio_core_outputs_lanedistributor_record6_we;
wire main_rtio_core_outputs_lanedistributor_record6_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record6_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record6_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record6_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record6_payload_data;
reg main_rtio_core_outputs_lanedistributor_record7_we;
wire main_rtio_core_outputs_lanedistributor_record7_writable;
wire [11:0] main_rtio_core_outputs_lanedistributor_record7_seqn;
wire [4:0] main_rtio_core_outputs_lanedistributor_record7_payload_channel;
reg [63:0] main_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
wire [7:0] main_rtio_core_outputs_lanedistributor_record7_payload_address;
wire [31:0] main_rtio_core_outputs_lanedistributor_record7_payload_data;
wire main_rtio_core_outputs_lanedistributor_o_status_wait;
reg main_rtio_core_outputs_lanedistributor_o_status_underflow = 1'd0;
reg [2:0] main_rtio_core_outputs_lanedistributor_current_lane = 3'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_coarse_timestamp = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 = 61'd0;
reg [60:0] main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 = 61'd0;
reg [11:0] main_rtio_core_outputs_lanedistributor_seqn = 12'd0;
wire [60:0] main_rtio_core_outputs_lanedistributor_coarse_timestamp;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_min_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp = 62'sd0;
reg signed [61:0] main_rtio_core_outputs_lanedistributor_last_minus_timestamp = 62'sd0;
wire [2:0] main_rtio_core_outputs_lanedistributor_current_lane_plus_one;
reg main_rtio_core_outputs_lanedistributor_quash = 1'd0;
wire [4:0] main_rtio_core_outputs_lanedistributor_adr;
wire [13:0] main_rtio_core_outputs_lanedistributor_dat_r;
wire signed [13:0] main_rtio_core_outputs_lanedistributor_compensation;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_last;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min;
wire main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min;
reg main_rtio_core_outputs_lanedistributor_force_laneB = 1'd0;
reg main_rtio_core_outputs_lanedistributor_use_laneB;
reg [2:0] main_rtio_core_outputs_lanedistributor_use_lanen;
reg main_rtio_core_outputs_lanedistributor_do_write;
reg main_rtio_core_outputs_lanedistributor_do_underflow;
reg main_rtio_core_outputs_lanedistributor_do_sequence_error;
wire [63:0] main_rtio_core_outputs_lanedistributor_compensated_timestamp;
wire main_rtio_core_outputs_lanedistributor_current_lane_writable;
reg main_rtio_core_outputs_lanedistributor_current_lane_writable_r = 1'd1;
wire main_rtio_core_outputs_record0_we;
wire main_rtio_core_outputs_record0_writable;
wire [11:0] main_rtio_core_outputs_record0_seqn0;
wire [4:0] main_rtio_core_outputs_record0_payload_channel0;
wire [63:0] main_rtio_core_outputs_record0_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record0_payload_address0;
wire [31:0] main_rtio_core_outputs_record0_payload_data0;
wire main_rtio_core_outputs_record1_we;
wire main_rtio_core_outputs_record1_writable;
wire [11:0] main_rtio_core_outputs_record1_seqn0;
wire [4:0] main_rtio_core_outputs_record1_payload_channel0;
wire [63:0] main_rtio_core_outputs_record1_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record1_payload_address0;
wire [31:0] main_rtio_core_outputs_record1_payload_data0;
wire main_rtio_core_outputs_record2_we;
wire main_rtio_core_outputs_record2_writable;
wire [11:0] main_rtio_core_outputs_record2_seqn0;
wire [4:0] main_rtio_core_outputs_record2_payload_channel0;
wire [63:0] main_rtio_core_outputs_record2_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record2_payload_address0;
wire [31:0] main_rtio_core_outputs_record2_payload_data0;
wire main_rtio_core_outputs_record3_we;
wire main_rtio_core_outputs_record3_writable;
wire [11:0] main_rtio_core_outputs_record3_seqn0;
wire [4:0] main_rtio_core_outputs_record3_payload_channel0;
wire [63:0] main_rtio_core_outputs_record3_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record3_payload_address0;
wire [31:0] main_rtio_core_outputs_record3_payload_data0;
wire main_rtio_core_outputs_record4_we;
wire main_rtio_core_outputs_record4_writable;
wire [11:0] main_rtio_core_outputs_record4_seqn0;
wire [4:0] main_rtio_core_outputs_record4_payload_channel0;
wire [63:0] main_rtio_core_outputs_record4_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record4_payload_address0;
wire [31:0] main_rtio_core_outputs_record4_payload_data0;
wire main_rtio_core_outputs_record5_we;
wire main_rtio_core_outputs_record5_writable;
wire [11:0] main_rtio_core_outputs_record5_seqn0;
wire [4:0] main_rtio_core_outputs_record5_payload_channel0;
wire [63:0] main_rtio_core_outputs_record5_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record5_payload_address0;
wire [31:0] main_rtio_core_outputs_record5_payload_data0;
wire main_rtio_core_outputs_record6_we;
wire main_rtio_core_outputs_record6_writable;
wire [11:0] main_rtio_core_outputs_record6_seqn0;
wire [4:0] main_rtio_core_outputs_record6_payload_channel0;
wire [63:0] main_rtio_core_outputs_record6_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record6_payload_address0;
wire [31:0] main_rtio_core_outputs_record6_payload_data0;
wire main_rtio_core_outputs_record7_we;
wire main_rtio_core_outputs_record7_writable;
wire [11:0] main_rtio_core_outputs_record7_seqn0;
wire [4:0] main_rtio_core_outputs_record7_payload_channel0;
wire [63:0] main_rtio_core_outputs_record7_payload_timestamp0;
wire [7:0] main_rtio_core_outputs_record7_payload_address0;
wire [31:0] main_rtio_core_outputs_record7_payload_data0;
wire main_rtio_core_outputs_record0_re;
wire main_rtio_core_outputs_record0_readable;
wire [11:0] main_rtio_core_outputs_record0_seqn1;
wire [4:0] main_rtio_core_outputs_record0_payload_channel1;
wire [63:0] main_rtio_core_outputs_record0_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record0_payload_address1;
wire [31:0] main_rtio_core_outputs_record0_payload_data1;
wire main_rtio_core_outputs_record1_re;
wire main_rtio_core_outputs_record1_readable;
wire [11:0] main_rtio_core_outputs_record1_seqn1;
wire [4:0] main_rtio_core_outputs_record1_payload_channel1;
wire [63:0] main_rtio_core_outputs_record1_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record1_payload_address1;
wire [31:0] main_rtio_core_outputs_record1_payload_data1;
wire main_rtio_core_outputs_record2_re;
wire main_rtio_core_outputs_record2_readable;
wire [11:0] main_rtio_core_outputs_record2_seqn1;
wire [4:0] main_rtio_core_outputs_record2_payload_channel1;
wire [63:0] main_rtio_core_outputs_record2_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record2_payload_address1;
wire [31:0] main_rtio_core_outputs_record2_payload_data1;
wire main_rtio_core_outputs_record3_re;
wire main_rtio_core_outputs_record3_readable;
wire [11:0] main_rtio_core_outputs_record3_seqn1;
wire [4:0] main_rtio_core_outputs_record3_payload_channel1;
wire [63:0] main_rtio_core_outputs_record3_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record3_payload_address1;
wire [31:0] main_rtio_core_outputs_record3_payload_data1;
wire main_rtio_core_outputs_record4_re;
wire main_rtio_core_outputs_record4_readable;
wire [11:0] main_rtio_core_outputs_record4_seqn1;
wire [4:0] main_rtio_core_outputs_record4_payload_channel1;
wire [63:0] main_rtio_core_outputs_record4_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record4_payload_address1;
wire [31:0] main_rtio_core_outputs_record4_payload_data1;
wire main_rtio_core_outputs_record5_re;
wire main_rtio_core_outputs_record5_readable;
wire [11:0] main_rtio_core_outputs_record5_seqn1;
wire [4:0] main_rtio_core_outputs_record5_payload_channel1;
wire [63:0] main_rtio_core_outputs_record5_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record5_payload_address1;
wire [31:0] main_rtio_core_outputs_record5_payload_data1;
wire main_rtio_core_outputs_record6_re;
wire main_rtio_core_outputs_record6_readable;
wire [11:0] main_rtio_core_outputs_record6_seqn1;
wire [4:0] main_rtio_core_outputs_record6_payload_channel1;
wire [63:0] main_rtio_core_outputs_record6_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record6_payload_address1;
wire [31:0] main_rtio_core_outputs_record6_payload_data1;
wire main_rtio_core_outputs_record7_re;
wire main_rtio_core_outputs_record7_readable;
wire [11:0] main_rtio_core_outputs_record7_seqn1;
wire [4:0] main_rtio_core_outputs_record7_payload_channel1;
wire [63:0] main_rtio_core_outputs_record7_payload_timestamp1;
wire [7:0] main_rtio_core_outputs_record7_payload_address1;
wire [31:0] main_rtio_core_outputs_record7_payload_data1;
wire main_rtio_core_outputs_asyncfifobuffered0_re;
reg main_rtio_core_outputs_asyncfifobuffered0_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered0_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re;
wire main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
wire main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered0_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered1_re;
reg main_rtio_core_outputs_asyncfifobuffered1_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered1_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re;
wire main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
wire main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered1_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered2_re;
reg main_rtio_core_outputs_asyncfifobuffered2_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered2_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re;
wire main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
wire main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered2_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered3_re;
reg main_rtio_core_outputs_asyncfifobuffered3_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered3_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re;
wire main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
wire main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered3_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered4_re;
reg main_rtio_core_outputs_asyncfifobuffered4_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered4_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re;
wire main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
wire main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered4_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered5_re;
reg main_rtio_core_outputs_asyncfifobuffered5_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered5_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re;
wire main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
wire main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered5_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered6_re;
reg main_rtio_core_outputs_asyncfifobuffered6_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered6_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re;
wire main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
wire main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered6_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered7_re;
reg main_rtio_core_outputs_asyncfifobuffered7_readable = 1'd0;
reg [120:0] main_rtio_core_outputs_asyncfifobuffered7_dout = 121'd0;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re;
wire main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
wire main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
wire main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q = 8'd0;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary = 8'd0;
reg [7:0] main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain;
wire [7:0] main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r;
wire main_rtio_core_outputs_asyncfifobuffered7_wrport_we;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
wire [6:0] main_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
wire [120:0] main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;
wire main_rtio_core_outputs_gates_record0_re;
wire main_rtio_core_outputs_gates_record0_readable;
wire [11:0] main_rtio_core_outputs_gates_record0_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record0_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record0_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record0_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record0_payload_data0;
wire main_rtio_core_outputs_gates_record1_re;
wire main_rtio_core_outputs_gates_record1_readable;
wire [11:0] main_rtio_core_outputs_gates_record1_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record1_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record1_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record1_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record1_payload_data0;
wire main_rtio_core_outputs_gates_record2_re;
wire main_rtio_core_outputs_gates_record2_readable;
wire [11:0] main_rtio_core_outputs_gates_record2_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record2_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record2_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record2_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record2_payload_data0;
wire main_rtio_core_outputs_gates_record3_re;
wire main_rtio_core_outputs_gates_record3_readable;
wire [11:0] main_rtio_core_outputs_gates_record3_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record3_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record3_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record3_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record3_payload_data0;
wire main_rtio_core_outputs_gates_record4_re;
wire main_rtio_core_outputs_gates_record4_readable;
wire [11:0] main_rtio_core_outputs_gates_record4_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record4_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record4_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record4_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record4_payload_data0;
wire main_rtio_core_outputs_gates_record5_re;
wire main_rtio_core_outputs_gates_record5_readable;
wire [11:0] main_rtio_core_outputs_gates_record5_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record5_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record5_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record5_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record5_payload_data0;
wire main_rtio_core_outputs_gates_record6_re;
wire main_rtio_core_outputs_gates_record6_readable;
wire [11:0] main_rtio_core_outputs_gates_record6_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record6_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record6_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record6_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record6_payload_data0;
wire main_rtio_core_outputs_gates_record7_re;
wire main_rtio_core_outputs_gates_record7_readable;
wire [11:0] main_rtio_core_outputs_gates_record7_seqn0;
wire [4:0] main_rtio_core_outputs_gates_record7_payload_channel0;
wire [63:0] main_rtio_core_outputs_gates_record7_payload_timestamp;
wire [7:0] main_rtio_core_outputs_gates_record7_payload_address0;
wire [31:0] main_rtio_core_outputs_gates_record7_payload_data0;
reg main_rtio_core_outputs_gates_record0_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record0_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record0_replace_occured;
wire main_rtio_core_outputs_gates_record0_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record0_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record0_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record0_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record0_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record1_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record1_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record1_replace_occured;
wire main_rtio_core_outputs_gates_record1_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record1_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record1_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record1_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record1_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record2_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record2_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record2_replace_occured;
wire main_rtio_core_outputs_gates_record2_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record2_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record2_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record2_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record2_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record3_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record3_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record3_replace_occured;
wire main_rtio_core_outputs_gates_record3_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record3_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record3_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record3_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record3_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record4_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record4_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record4_replace_occured;
wire main_rtio_core_outputs_gates_record4_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record4_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record4_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record4_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record4_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record5_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record5_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record5_replace_occured;
wire main_rtio_core_outputs_gates_record5_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record5_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record5_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record5_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record5_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record6_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record6_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record6_replace_occured;
wire main_rtio_core_outputs_gates_record6_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record6_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record6_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record6_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record6_payload_data1 = 32'd0;
reg main_rtio_core_outputs_gates_record7_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_gates_record7_seqn1 = 12'd0;
wire main_rtio_core_outputs_gates_record7_replace_occured;
wire main_rtio_core_outputs_gates_record7_nondata_replace_occured;
reg [4:0] main_rtio_core_outputs_gates_record7_payload_channel1 = 5'd0;
reg [2:0] main_rtio_core_outputs_gates_record7_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_gates_record7_payload_address1 = 8'd0;
reg [31:0] main_rtio_core_outputs_gates_record7_payload_data1 = 32'd0;
wire [60:0] main_rtio_core_outputs_gates_coarse_timestamp;
reg main_rtio_core_outputs_collision = 1'd0;
reg [4:0] main_rtio_core_outputs_collision_channel = 5'd0;
reg main_rtio_core_outputs_busy = 1'd0;
reg [4:0] main_rtio_core_outputs_busy_channel = 5'd0;
wire main_rtio_core_outputs_record0_valid0;
wire [11:0] main_rtio_core_outputs_record0_seqn2;
wire main_rtio_core_outputs_record0_replace_occured;
wire main_rtio_core_outputs_record0_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record0_payload_channel2;
wire [2:0] main_rtio_core_outputs_record0_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record0_payload_address2;
wire [31:0] main_rtio_core_outputs_record0_payload_data2;
wire main_rtio_core_outputs_record1_valid0;
wire [11:0] main_rtio_core_outputs_record1_seqn2;
wire main_rtio_core_outputs_record1_replace_occured;
wire main_rtio_core_outputs_record1_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record1_payload_channel2;
wire [2:0] main_rtio_core_outputs_record1_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record1_payload_address2;
wire [31:0] main_rtio_core_outputs_record1_payload_data2;
wire main_rtio_core_outputs_record2_valid0;
wire [11:0] main_rtio_core_outputs_record2_seqn2;
wire main_rtio_core_outputs_record2_replace_occured;
wire main_rtio_core_outputs_record2_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record2_payload_channel2;
wire [2:0] main_rtio_core_outputs_record2_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record2_payload_address2;
wire [31:0] main_rtio_core_outputs_record2_payload_data2;
wire main_rtio_core_outputs_record3_valid0;
wire [11:0] main_rtio_core_outputs_record3_seqn2;
wire main_rtio_core_outputs_record3_replace_occured;
wire main_rtio_core_outputs_record3_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record3_payload_channel2;
wire [2:0] main_rtio_core_outputs_record3_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record3_payload_address2;
wire [31:0] main_rtio_core_outputs_record3_payload_data2;
wire main_rtio_core_outputs_record4_valid0;
wire [11:0] main_rtio_core_outputs_record4_seqn2;
wire main_rtio_core_outputs_record4_replace_occured;
wire main_rtio_core_outputs_record4_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record4_payload_channel2;
wire [2:0] main_rtio_core_outputs_record4_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record4_payload_address2;
wire [31:0] main_rtio_core_outputs_record4_payload_data2;
wire main_rtio_core_outputs_record5_valid0;
wire [11:0] main_rtio_core_outputs_record5_seqn2;
wire main_rtio_core_outputs_record5_replace_occured;
wire main_rtio_core_outputs_record5_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record5_payload_channel2;
wire [2:0] main_rtio_core_outputs_record5_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record5_payload_address2;
wire [31:0] main_rtio_core_outputs_record5_payload_data2;
wire main_rtio_core_outputs_record6_valid0;
wire [11:0] main_rtio_core_outputs_record6_seqn2;
wire main_rtio_core_outputs_record6_replace_occured;
wire main_rtio_core_outputs_record6_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record6_payload_channel2;
wire [2:0] main_rtio_core_outputs_record6_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record6_payload_address2;
wire [31:0] main_rtio_core_outputs_record6_payload_data2;
wire main_rtio_core_outputs_record7_valid0;
wire [11:0] main_rtio_core_outputs_record7_seqn2;
wire main_rtio_core_outputs_record7_replace_occured;
wire main_rtio_core_outputs_record7_nondata_replace_occured;
wire [4:0] main_rtio_core_outputs_record7_payload_channel2;
wire [2:0] main_rtio_core_outputs_record7_payload_fine_ts0;
wire [7:0] main_rtio_core_outputs_record7_payload_address2;
wire [31:0] main_rtio_core_outputs_record7_payload_data2;
reg main_rtio_core_outputs_record0_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record0_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record0_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record0_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record0_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record0_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record0_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record0_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record1_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record1_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record1_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record1_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record1_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record1_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record1_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record1_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record2_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record2_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record2_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record2_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record2_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record2_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record2_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record2_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record3_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record3_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record3_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record3_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record3_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record3_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record3_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record3_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record4_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record4_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record4_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record4_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record4_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record4_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record4_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record4_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record5_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record5_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record5_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record5_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record5_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record5_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record5_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record5_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record6_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record6_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record6_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record6_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record6_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record6_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record6_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record6_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record7_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record7_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record7_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record7_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record7_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record7_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record7_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record7_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference0;
reg main_rtio_core_outputs_nondata_difference1;
reg main_rtio_core_outputs_nondata_difference2;
reg main_rtio_core_outputs_nondata_difference3;
reg main_rtio_core_outputs_record8_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record8_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record8_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record8_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record8_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record8_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record8_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record8_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record9_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record9_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record9_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record9_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record9_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record9_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record9_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record9_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record10_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record10_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record10_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record10_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record10_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record10_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record10_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record10_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record11_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record11_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record11_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record11_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record11_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record11_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record11_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record11_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record12_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record12_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record12_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record12_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record12_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record12_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record12_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record12_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record13_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record13_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record13_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record13_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record13_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record13_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record13_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record13_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record14_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record14_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record14_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record14_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record14_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record14_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record14_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record14_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record15_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record15_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record15_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record15_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record15_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record15_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record15_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record15_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference4;
reg main_rtio_core_outputs_nondata_difference5;
reg main_rtio_core_outputs_nondata_difference6;
reg main_rtio_core_outputs_nondata_difference7;
reg main_rtio_core_outputs_record16_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record16_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record16_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record16_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record16_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record16_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record16_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record16_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record17_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record17_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record17_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record17_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record17_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record17_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record17_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record17_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record18_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record18_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record18_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record18_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record18_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record18_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record18_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record18_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record19_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record19_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record19_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record19_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record19_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record19_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record19_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record19_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record20_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record20_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record20_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record20_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record20_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record20_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record20_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record20_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record21_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record21_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record21_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record21_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record21_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record21_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record21_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record21_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record22_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record22_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record22_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record22_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record22_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record22_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record22_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record22_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record23_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record23_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record23_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record23_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record23_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record23_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record23_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record23_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference8;
reg main_rtio_core_outputs_nondata_difference9;
reg main_rtio_core_outputs_record24_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record24_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record24_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record24_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record24_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record24_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record24_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record24_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record25_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record25_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record25_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record25_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record25_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record25_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record25_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record25_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record26_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record26_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record26_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record26_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record26_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record26_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record26_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record26_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record27_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record27_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record27_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record27_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record27_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record27_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record27_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record27_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record28_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record28_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record28_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record28_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record28_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record28_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record28_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record28_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record29_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record29_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record29_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record29_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record29_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record29_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record29_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record29_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record30_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record30_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record30_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record30_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record30_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record30_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record30_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record30_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record31_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record31_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record31_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record31_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record31_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record31_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record31_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record31_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference10;
reg main_rtio_core_outputs_nondata_difference11;
reg main_rtio_core_outputs_nondata_difference12;
reg main_rtio_core_outputs_nondata_difference13;
reg main_rtio_core_outputs_record32_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record32_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record32_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record32_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record32_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record32_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record32_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record32_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record33_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record33_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record33_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record33_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record33_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record33_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record33_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record33_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record34_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record34_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record34_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record34_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record34_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record34_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record34_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record34_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record35_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record35_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record35_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record35_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record35_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record35_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record35_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record35_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record36_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record36_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record36_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record36_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record36_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record36_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record36_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record36_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record37_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record37_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record37_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record37_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record37_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record37_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record37_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record37_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record38_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record38_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record38_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record38_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record38_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record38_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record38_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record38_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record39_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record39_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record39_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record39_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record39_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record39_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record39_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record39_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference14;
reg main_rtio_core_outputs_nondata_difference15;
reg main_rtio_core_outputs_record40_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record40_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record40_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record40_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record40_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record40_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record40_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record40_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record41_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record41_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record41_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record41_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record41_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record41_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record41_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record41_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record42_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record42_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record42_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record42_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record42_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record42_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record42_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record42_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record43_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record43_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record43_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record43_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record43_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record43_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record43_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record43_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record44_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record44_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record44_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record44_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record44_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record44_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record44_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record44_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record45_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record45_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record45_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record45_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record45_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record45_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record45_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record45_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record46_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record46_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record46_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record46_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record46_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record46_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record46_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record46_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_record47_rec_valid = 1'd0;
reg [11:0] main_rtio_core_outputs_record47_rec_seqn = 12'd0;
reg main_rtio_core_outputs_record47_rec_replace_occured = 1'd0;
reg main_rtio_core_outputs_record47_rec_nondata_replace_occured = 1'd0;
reg [4:0] main_rtio_core_outputs_record47_rec_payload_channel = 5'd0;
reg [2:0] main_rtio_core_outputs_record47_rec_payload_fine_ts = 3'd0;
reg [7:0] main_rtio_core_outputs_record47_rec_payload_address = 8'd0;
reg [31:0] main_rtio_core_outputs_record47_rec_payload_data = 32'd0;
reg main_rtio_core_outputs_nondata_difference16;
reg main_rtio_core_outputs_nondata_difference17;
reg main_rtio_core_outputs_nondata_difference18;
reg main_rtio_core_outputs_record0_valid1 = 1'd0;
wire main_rtio_core_outputs_record0_collision;
reg [4:0] main_rtio_core_outputs_record0_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record0_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record0_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record0_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record1_valid1 = 1'd0;
wire main_rtio_core_outputs_record1_collision;
reg [4:0] main_rtio_core_outputs_record1_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record1_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record1_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record1_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record2_valid1 = 1'd0;
wire main_rtio_core_outputs_record2_collision;
reg [4:0] main_rtio_core_outputs_record2_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record2_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record2_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record2_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record3_valid1 = 1'd0;
wire main_rtio_core_outputs_record3_collision;
reg [4:0] main_rtio_core_outputs_record3_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record3_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record3_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record3_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record4_valid1 = 1'd0;
wire main_rtio_core_outputs_record4_collision;
reg [4:0] main_rtio_core_outputs_record4_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record4_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record4_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record4_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record5_valid1 = 1'd0;
wire main_rtio_core_outputs_record5_collision;
reg [4:0] main_rtio_core_outputs_record5_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record5_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record5_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record5_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record6_valid1 = 1'd0;
wire main_rtio_core_outputs_record6_collision;
reg [4:0] main_rtio_core_outputs_record6_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record6_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record6_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record6_payload_data3 = 32'd0;
reg main_rtio_core_outputs_record7_valid1 = 1'd0;
wire main_rtio_core_outputs_record7_collision;
reg [4:0] main_rtio_core_outputs_record7_payload_channel3 = 5'd0;
reg [2:0] main_rtio_core_outputs_record7_payload_fine_ts1 = 3'd0;
reg [7:0] main_rtio_core_outputs_record7_payload_address3 = 8'd0;
reg [31:0] main_rtio_core_outputs_record7_payload_data3 = 32'd0;
reg main_rtio_core_outputs_replace_occured_r0 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r0 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory0_adr;
wire main_rtio_core_outputs_memory0_dat_r;
reg main_rtio_core_outputs_replace_occured_r1 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r1 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory1_adr;
wire main_rtio_core_outputs_memory1_dat_r;
reg main_rtio_core_outputs_replace_occured_r2 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r2 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory2_adr;
wire main_rtio_core_outputs_memory2_dat_r;
reg main_rtio_core_outputs_replace_occured_r3 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r3 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory3_adr;
wire main_rtio_core_outputs_memory3_dat_r;
reg main_rtio_core_outputs_replace_occured_r4 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r4 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory4_adr;
wire main_rtio_core_outputs_memory4_dat_r;
reg main_rtio_core_outputs_replace_occured_r5 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r5 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory5_adr;
wire main_rtio_core_outputs_memory5_dat_r;
reg main_rtio_core_outputs_replace_occured_r6 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r6 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory6_adr;
wire main_rtio_core_outputs_memory6_dat_r;
reg main_rtio_core_outputs_replace_occured_r7 = 1'd0;
reg main_rtio_core_outputs_nondata_replace_occured_r7 = 1'd0;
wire [4:0] main_rtio_core_outputs_memory7_adr;
wire main_rtio_core_outputs_memory7_dat_r;
wire main_rtio_core_outputs_selected0;
wire main_rtio_core_outputs_selected1;
wire main_rtio_core_outputs_selected2;
wire main_rtio_core_outputs_selected3;
wire main_rtio_core_outputs_selected4;
wire main_rtio_core_outputs_selected5;
wire main_rtio_core_outputs_selected6;
wire main_rtio_core_outputs_selected7;
wire main_rtio_core_outputs_selected8;
wire main_rtio_core_outputs_selected9;
wire main_rtio_core_outputs_selected10;
wire main_rtio_core_outputs_selected11;
wire main_rtio_core_outputs_selected12;
wire main_rtio_core_outputs_selected13;
wire main_rtio_core_outputs_selected14;
wire main_rtio_core_outputs_selected15;
wire main_rtio_core_outputs_selected16;
wire main_rtio_core_outputs_selected17;
wire main_rtio_core_outputs_selected18;
wire main_rtio_core_outputs_selected19;
wire main_rtio_core_outputs_selected20;
wire main_rtio_core_outputs_selected21;
wire main_rtio_core_outputs_selected22;
wire main_rtio_core_outputs_selected23;
wire main_rtio_core_outputs_selected24;
wire main_rtio_core_outputs_selected25;
wire main_rtio_core_outputs_selected26;
wire main_rtio_core_outputs_selected27;
wire main_rtio_core_outputs_selected28;
wire main_rtio_core_outputs_selected29;
wire main_rtio_core_outputs_selected30;
wire main_rtio_core_outputs_selected31;
wire main_rtio_core_outputs_selected32;
wire main_rtio_core_outputs_selected33;
wire main_rtio_core_outputs_selected34;
wire main_rtio_core_outputs_selected35;
wire main_rtio_core_outputs_selected36;
wire main_rtio_core_outputs_selected37;
wire main_rtio_core_outputs_selected38;
wire main_rtio_core_outputs_selected39;
wire main_rtio_core_outputs_selected40;
wire main_rtio_core_outputs_selected41;
wire main_rtio_core_outputs_selected42;
wire main_rtio_core_outputs_selected43;
wire main_rtio_core_outputs_selected44;
wire main_rtio_core_outputs_selected45;
wire main_rtio_core_outputs_selected46;
wire main_rtio_core_outputs_selected47;
wire main_rtio_core_outputs_selected48;
wire main_rtio_core_outputs_selected49;
wire main_rtio_core_outputs_selected50;
wire main_rtio_core_outputs_selected51;
wire main_rtio_core_outputs_selected52;
wire main_rtio_core_outputs_selected53;
wire main_rtio_core_outputs_selected54;
wire main_rtio_core_outputs_selected55;
wire main_rtio_core_outputs_selected56;
wire main_rtio_core_outputs_selected57;
wire main_rtio_core_outputs_selected58;
wire main_rtio_core_outputs_selected59;
wire main_rtio_core_outputs_selected60;
wire main_rtio_core_outputs_selected61;
wire main_rtio_core_outputs_selected62;
wire main_rtio_core_outputs_selected63;
wire main_rtio_core_outputs_selected64;
wire main_rtio_core_outputs_selected65;
wire main_rtio_core_outputs_selected66;
wire main_rtio_core_outputs_selected67;
wire main_rtio_core_outputs_selected68;
wire main_rtio_core_outputs_selected69;
wire main_rtio_core_outputs_selected70;
wire main_rtio_core_outputs_selected71;
wire main_rtio_core_outputs_selected72;
wire main_rtio_core_outputs_selected73;
wire main_rtio_core_outputs_selected74;
wire main_rtio_core_outputs_selected75;
wire main_rtio_core_outputs_selected76;
wire main_rtio_core_outputs_selected77;
wire main_rtio_core_outputs_selected78;
wire main_rtio_core_outputs_selected79;
wire main_rtio_core_outputs_selected80;
wire main_rtio_core_outputs_selected81;
wire main_rtio_core_outputs_selected82;
wire main_rtio_core_outputs_selected83;
wire main_rtio_core_outputs_selected84;
wire main_rtio_core_outputs_selected85;
wire main_rtio_core_outputs_selected86;
wire main_rtio_core_outputs_selected87;
wire main_rtio_core_outputs_selected88;
wire main_rtio_core_outputs_selected89;
wire main_rtio_core_outputs_selected90;
wire main_rtio_core_outputs_selected91;
wire main_rtio_core_outputs_selected92;
wire main_rtio_core_outputs_selected93;
wire main_rtio_core_outputs_selected94;
wire main_rtio_core_outputs_selected95;
wire main_rtio_core_outputs_selected96;
wire main_rtio_core_outputs_selected97;
wire main_rtio_core_outputs_selected98;
wire main_rtio_core_outputs_selected99;
wire main_rtio_core_outputs_selected100;
wire main_rtio_core_outputs_selected101;
wire main_rtio_core_outputs_selected102;
wire main_rtio_core_outputs_selected103;
wire main_rtio_core_outputs_selected104;
wire main_rtio_core_outputs_selected105;
wire main_rtio_core_outputs_selected106;
wire main_rtio_core_outputs_selected107;
wire main_rtio_core_outputs_selected108;
wire main_rtio_core_outputs_selected109;
wire main_rtio_core_outputs_selected110;
wire main_rtio_core_outputs_selected111;
wire main_rtio_core_outputs_selected112;
wire main_rtio_core_outputs_selected113;
wire main_rtio_core_outputs_selected114;
wire main_rtio_core_outputs_selected115;
wire main_rtio_core_outputs_selected116;
wire main_rtio_core_outputs_selected117;
wire main_rtio_core_outputs_selected118;
wire main_rtio_core_outputs_selected119;
wire main_rtio_core_outputs_selected120;
wire main_rtio_core_outputs_selected121;
wire main_rtio_core_outputs_selected122;
wire main_rtio_core_outputs_selected123;
wire main_rtio_core_outputs_selected124;
wire main_rtio_core_outputs_selected125;
wire main_rtio_core_outputs_selected126;
wire main_rtio_core_outputs_selected127;
wire main_rtio_core_outputs_selected128;
wire main_rtio_core_outputs_selected129;
wire main_rtio_core_outputs_selected130;
wire main_rtio_core_outputs_selected131;
wire main_rtio_core_outputs_selected132;
wire main_rtio_core_outputs_selected133;
wire main_rtio_core_outputs_selected134;
wire main_rtio_core_outputs_selected135;
wire main_rtio_core_outputs_selected136;
wire main_rtio_core_outputs_selected137;
wire main_rtio_core_outputs_selected138;
wire main_rtio_core_outputs_selected139;
wire main_rtio_core_outputs_selected140;
wire main_rtio_core_outputs_selected141;
wire main_rtio_core_outputs_selected142;
wire main_rtio_core_outputs_selected143;
wire main_rtio_core_outputs_selected144;
wire main_rtio_core_outputs_selected145;
wire main_rtio_core_outputs_selected146;
wire main_rtio_core_outputs_selected147;
wire main_rtio_core_outputs_selected148;
wire main_rtio_core_outputs_selected149;
wire main_rtio_core_outputs_selected150;
wire main_rtio_core_outputs_selected151;
wire main_rtio_core_outputs_selected152;
wire main_rtio_core_outputs_selected153;
wire main_rtio_core_outputs_selected154;
wire main_rtio_core_outputs_selected155;
wire main_rtio_core_outputs_selected156;
wire main_rtio_core_outputs_selected157;
wire main_rtio_core_outputs_selected158;
wire main_rtio_core_outputs_selected159;
wire main_rtio_core_outputs_selected160;
wire main_rtio_core_outputs_selected161;
wire main_rtio_core_outputs_selected162;
wire main_rtio_core_outputs_selected163;
wire main_rtio_core_outputs_selected164;
wire main_rtio_core_outputs_selected165;
wire main_rtio_core_outputs_selected166;
wire main_rtio_core_outputs_selected167;
wire main_rtio_core_outputs_selected168;
wire main_rtio_core_outputs_selected169;
wire main_rtio_core_outputs_selected170;
wire main_rtio_core_outputs_selected171;
wire main_rtio_core_outputs_selected172;
wire main_rtio_core_outputs_selected173;
wire main_rtio_core_outputs_selected174;
wire main_rtio_core_outputs_selected175;
wire main_rtio_core_outputs_selected176;
wire main_rtio_core_outputs_selected177;
wire main_rtio_core_outputs_selected178;
wire main_rtio_core_outputs_selected179;
wire main_rtio_core_outputs_selected180;
wire main_rtio_core_outputs_selected181;
wire main_rtio_core_outputs_selected182;
wire main_rtio_core_outputs_selected183;
wire main_rtio_core_outputs_selected184;
wire main_rtio_core_outputs_selected185;
wire main_rtio_core_outputs_selected186;
wire main_rtio_core_outputs_selected187;
wire main_rtio_core_outputs_selected188;
wire main_rtio_core_outputs_selected189;
wire main_rtio_core_outputs_selected190;
wire main_rtio_core_outputs_selected191;
wire main_rtio_core_outputs_selected192;
wire main_rtio_core_outputs_selected193;
wire main_rtio_core_outputs_selected194;
wire main_rtio_core_outputs_selected195;
wire main_rtio_core_outputs_selected196;
wire main_rtio_core_outputs_selected197;
wire main_rtio_core_outputs_selected198;
wire main_rtio_core_outputs_selected199;
wire main_rtio_core_outputs_selected200;
wire main_rtio_core_outputs_selected201;
wire main_rtio_core_outputs_selected202;
wire main_rtio_core_outputs_selected203;
wire main_rtio_core_outputs_selected204;
wire main_rtio_core_outputs_selected205;
wire main_rtio_core_outputs_selected206;
wire main_rtio_core_outputs_selected207;
wire main_rtio_core_outputs_selected208;
wire main_rtio_core_outputs_selected209;
wire main_rtio_core_outputs_selected210;
wire main_rtio_core_outputs_selected211;
wire main_rtio_core_outputs_selected212;
wire main_rtio_core_outputs_selected213;
wire main_rtio_core_outputs_selected214;
wire main_rtio_core_outputs_selected215;
wire main_rtio_core_outputs_selected216;
wire main_rtio_core_outputs_selected217;
wire main_rtio_core_outputs_selected218;
wire main_rtio_core_outputs_selected219;
wire main_rtio_core_outputs_selected220;
wire main_rtio_core_outputs_selected221;
wire main_rtio_core_outputs_selected222;
wire main_rtio_core_outputs_selected223;
wire main_rtio_core_outputs_selected224;
wire main_rtio_core_outputs_selected225;
wire main_rtio_core_outputs_selected226;
wire main_rtio_core_outputs_selected227;
wire main_rtio_core_outputs_selected228;
wire main_rtio_core_outputs_selected229;
wire main_rtio_core_outputs_selected230;
wire main_rtio_core_outputs_selected231;
reg main_rtio_core_outputs_stb_r0 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r0 = 5'd0;
reg main_rtio_core_outputs_stb_r1 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r1 = 5'd0;
reg main_rtio_core_outputs_stb_r2 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r2 = 5'd0;
reg main_rtio_core_outputs_stb_r3 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r3 = 5'd0;
reg main_rtio_core_outputs_stb_r4 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r4 = 5'd0;
reg main_rtio_core_outputs_stb_r5 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r5 = 5'd0;
reg main_rtio_core_outputs_stb_r6 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r6 = 5'd0;
reg main_rtio_core_outputs_stb_r7 = 1'd0;
reg [4:0] main_rtio_core_outputs_channel_r7 = 5'd0;
reg main_rtio_core_inputs_i_ack = 1'd0;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_we;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_re;
wire main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
wire [64:0] main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
wire main_rtio_core_inputs_asyncfifo0_graycounter0_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
wire main_rtio_core_inputs_asyncfifo0_graycounter1_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo0_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo0_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo0_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo0_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo0_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo0_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo0_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo0_rdport_dat_r;
wire main_rtio_core_inputs_record0_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record0_fifo_in_timestamp;
wire main_rtio_core_inputs_record0_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record0_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io0;
wire main_rtio_core_inputs_blindtransfer0_i;
wire main_rtio_core_inputs_blindtransfer0_o;
wire main_rtio_core_inputs_blindtransfer0_ps_i;
wire main_rtio_core_inputs_blindtransfer0_ps_o;
reg main_rtio_core_inputs_blindtransfer0_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer0_blind = 1'd0;
wire main_rtio_core_inputs_selected0;
reg main_rtio_core_inputs_overflow0 = 1'd0;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_we;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_re;
wire main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
wire [64:0] main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
wire main_rtio_core_inputs_asyncfifo1_graycounter2_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
wire main_rtio_core_inputs_asyncfifo1_graycounter3_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo1_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo1_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo1_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo1_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo1_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo1_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo1_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo1_rdport_dat_r;
wire main_rtio_core_inputs_record1_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record1_fifo_in_timestamp;
wire main_rtio_core_inputs_record1_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record1_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io1;
wire main_rtio_core_inputs_blindtransfer1_i;
wire main_rtio_core_inputs_blindtransfer1_o;
wire main_rtio_core_inputs_blindtransfer1_ps_i;
wire main_rtio_core_inputs_blindtransfer1_ps_o;
reg main_rtio_core_inputs_blindtransfer1_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer1_blind = 1'd0;
wire main_rtio_core_inputs_selected1;
reg main_rtio_core_inputs_overflow1 = 1'd0;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_we;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_re;
wire main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
wire [64:0] main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
wire main_rtio_core_inputs_asyncfifo2_graycounter4_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
wire main_rtio_core_inputs_asyncfifo2_graycounter5_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo2_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo2_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo2_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo2_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo2_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo2_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo2_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo2_rdport_dat_r;
wire main_rtio_core_inputs_record2_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record2_fifo_in_timestamp;
wire main_rtio_core_inputs_record2_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record2_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io2;
wire main_rtio_core_inputs_blindtransfer2_i;
wire main_rtio_core_inputs_blindtransfer2_o;
wire main_rtio_core_inputs_blindtransfer2_ps_i;
wire main_rtio_core_inputs_blindtransfer2_ps_o;
reg main_rtio_core_inputs_blindtransfer2_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer2_blind = 1'd0;
wire main_rtio_core_inputs_selected2;
reg main_rtio_core_inputs_overflow2 = 1'd0;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_we;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_re;
wire main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
wire [64:0] main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
wire main_rtio_core_inputs_asyncfifo3_graycounter6_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
wire main_rtio_core_inputs_asyncfifo3_graycounter7_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo3_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo3_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo3_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo3_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo3_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo3_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo3_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo3_rdport_dat_r;
wire main_rtio_core_inputs_record3_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record3_fifo_in_timestamp;
wire main_rtio_core_inputs_record3_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record3_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io3;
wire main_rtio_core_inputs_blindtransfer3_i;
wire main_rtio_core_inputs_blindtransfer3_o;
wire main_rtio_core_inputs_blindtransfer3_ps_i;
wire main_rtio_core_inputs_blindtransfer3_ps_o;
reg main_rtio_core_inputs_blindtransfer3_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer3_blind = 1'd0;
wire main_rtio_core_inputs_selected3;
reg main_rtio_core_inputs_overflow3 = 1'd0;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_we;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_re;
wire main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
wire [64:0] main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
wire main_rtio_core_inputs_asyncfifo4_graycounter8_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
wire main_rtio_core_inputs_asyncfifo4_graycounter9_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo4_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo4_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo4_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo4_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo4_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo4_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo4_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo4_rdport_dat_r;
wire main_rtio_core_inputs_record4_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record4_fifo_in_timestamp;
wire main_rtio_core_inputs_record4_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record4_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io4;
wire main_rtio_core_inputs_blindtransfer4_i;
wire main_rtio_core_inputs_blindtransfer4_o;
wire main_rtio_core_inputs_blindtransfer4_ps_i;
wire main_rtio_core_inputs_blindtransfer4_ps_o;
reg main_rtio_core_inputs_blindtransfer4_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer4_blind = 1'd0;
wire main_rtio_core_inputs_selected4;
reg main_rtio_core_inputs_overflow4 = 1'd0;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_we;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_re;
wire main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
wire [64:0] main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
wire main_rtio_core_inputs_asyncfifo5_graycounter10_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
wire main_rtio_core_inputs_asyncfifo5_graycounter11_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo5_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo5_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo5_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo5_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo5_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo5_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo5_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo5_rdport_dat_r;
wire main_rtio_core_inputs_record5_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record5_fifo_in_timestamp;
wire main_rtio_core_inputs_record5_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record5_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io5;
wire main_rtio_core_inputs_blindtransfer5_i;
wire main_rtio_core_inputs_blindtransfer5_o;
wire main_rtio_core_inputs_blindtransfer5_ps_i;
wire main_rtio_core_inputs_blindtransfer5_ps_o;
reg main_rtio_core_inputs_blindtransfer5_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer5_blind = 1'd0;
wire main_rtio_core_inputs_selected5;
reg main_rtio_core_inputs_overflow5 = 1'd0;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_we;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_re;
wire main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable;
wire [64:0] main_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
wire [64:0] main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
wire main_rtio_core_inputs_asyncfifo6_graycounter12_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
wire main_rtio_core_inputs_asyncfifo6_graycounter13_ce;
(* dont_touch = "true" *) reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q = 10'd0;
wire [9:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary = 10'd0;
reg [9:0] main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
wire [9:0] main_rtio_core_inputs_asyncfifo6_produce_rdomain;
wire [9:0] main_rtio_core_inputs_asyncfifo6_consume_wdomain;
wire [8:0] main_rtio_core_inputs_asyncfifo6_wrport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo6_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo6_wrport_we;
wire [64:0] main_rtio_core_inputs_asyncfifo6_wrport_dat_w;
wire [8:0] main_rtio_core_inputs_asyncfifo6_rdport_adr;
wire [64:0] main_rtio_core_inputs_asyncfifo6_rdport_dat_r;
wire main_rtio_core_inputs_record6_fifo_in_data;
wire [63:0] main_rtio_core_inputs_record6_fifo_in_timestamp;
wire main_rtio_core_inputs_record6_fifo_out_data;
wire [63:0] main_rtio_core_inputs_record6_fifo_out_timestamp;
wire main_rtio_core_inputs_overflow_io6;
wire main_rtio_core_inputs_blindtransfer6_i;
wire main_rtio_core_inputs_blindtransfer6_o;
wire main_rtio_core_inputs_blindtransfer6_ps_i;
wire main_rtio_core_inputs_blindtransfer6_ps_o;
reg main_rtio_core_inputs_blindtransfer6_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer6_blind = 1'd0;
wire main_rtio_core_inputs_selected6;
reg main_rtio_core_inputs_overflow6 = 1'd0;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_we;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_re;
wire main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo7_asyncfifo7_din;
wire [31:0] main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout;
wire main_rtio_core_inputs_asyncfifo7_graycounter14_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary;
wire main_rtio_core_inputs_asyncfifo7_graycounter15_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary;
wire [2:0] main_rtio_core_inputs_asyncfifo7_produce_rdomain;
wire [2:0] main_rtio_core_inputs_asyncfifo7_consume_wdomain;
wire [1:0] main_rtio_core_inputs_asyncfifo7_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo7_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo7_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo7_wrport_dat_w;
wire [1:0] main_rtio_core_inputs_asyncfifo7_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo7_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record7_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record7_fifo_out_data;
wire main_rtio_core_inputs_overflow_io7;
wire main_rtio_core_inputs_blindtransfer7_i;
wire main_rtio_core_inputs_blindtransfer7_o;
wire main_rtio_core_inputs_blindtransfer7_ps_i;
wire main_rtio_core_inputs_blindtransfer7_ps_o;
reg main_rtio_core_inputs_blindtransfer7_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer7_blind = 1'd0;
wire main_rtio_core_inputs_selected7;
reg main_rtio_core_inputs_overflow7 = 1'd0;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_we;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_re;
wire main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo8_asyncfifo8_din;
wire [31:0] main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout;
wire main_rtio_core_inputs_asyncfifo8_graycounter16_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary;
wire main_rtio_core_inputs_asyncfifo8_graycounter17_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary;
wire [7:0] main_rtio_core_inputs_asyncfifo8_produce_rdomain;
wire [7:0] main_rtio_core_inputs_asyncfifo8_consume_wdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo8_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo8_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo8_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo8_wrport_dat_w;
wire [6:0] main_rtio_core_inputs_asyncfifo8_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo8_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record8_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record8_fifo_out_data;
wire main_rtio_core_inputs_overflow_io8;
wire main_rtio_core_inputs_blindtransfer8_i;
wire main_rtio_core_inputs_blindtransfer8_o;
wire main_rtio_core_inputs_blindtransfer8_ps_i;
wire main_rtio_core_inputs_blindtransfer8_ps_o;
reg main_rtio_core_inputs_blindtransfer8_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer8_blind = 1'd0;
wire main_rtio_core_inputs_selected8;
reg main_rtio_core_inputs_overflow8 = 1'd0;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_we;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_re;
wire main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo9_asyncfifo9_din;
wire [31:0] main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout;
wire main_rtio_core_inputs_asyncfifo9_graycounter18_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary;
wire main_rtio_core_inputs_asyncfifo9_graycounter19_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary;
wire [7:0] main_rtio_core_inputs_asyncfifo9_produce_rdomain;
wire [7:0] main_rtio_core_inputs_asyncfifo9_consume_wdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo9_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo9_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo9_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo9_wrport_dat_w;
wire [6:0] main_rtio_core_inputs_asyncfifo9_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo9_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record9_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record9_fifo_out_data;
wire main_rtio_core_inputs_overflow_io9;
wire main_rtio_core_inputs_blindtransfer9_i;
wire main_rtio_core_inputs_blindtransfer9_o;
wire main_rtio_core_inputs_blindtransfer9_ps_i;
wire main_rtio_core_inputs_blindtransfer9_ps_o;
reg main_rtio_core_inputs_blindtransfer9_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer9_blind = 1'd0;
wire main_rtio_core_inputs_selected9;
reg main_rtio_core_inputs_overflow9 = 1'd0;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_we;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_re;
wire main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo10_asyncfifo10_din;
wire [31:0] main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout;
wire main_rtio_core_inputs_asyncfifo10_graycounter20_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary;
wire main_rtio_core_inputs_asyncfifo10_graycounter21_ce;
(* dont_touch = "true" *) reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q = 8'd0;
wire [7:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_next;
reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary = 8'd0;
reg [7:0] main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary;
wire [7:0] main_rtio_core_inputs_asyncfifo10_produce_rdomain;
wire [7:0] main_rtio_core_inputs_asyncfifo10_consume_wdomain;
wire [6:0] main_rtio_core_inputs_asyncfifo10_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo10_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo10_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo10_wrport_dat_w;
wire [6:0] main_rtio_core_inputs_asyncfifo10_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo10_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record10_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record10_fifo_out_data;
wire main_rtio_core_inputs_overflow_io10;
wire main_rtio_core_inputs_blindtransfer10_i;
wire main_rtio_core_inputs_blindtransfer10_o;
wire main_rtio_core_inputs_blindtransfer10_ps_i;
wire main_rtio_core_inputs_blindtransfer10_ps_o;
reg main_rtio_core_inputs_blindtransfer10_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer10_blind = 1'd0;
wire main_rtio_core_inputs_selected10;
reg main_rtio_core_inputs_overflow10 = 1'd0;
wire main_rtio_core_inputs_asyncfifo11_asyncfifo11_we;
wire main_rtio_core_inputs_asyncfifo11_asyncfifo11_writable;
wire main_rtio_core_inputs_asyncfifo11_asyncfifo11_re;
wire main_rtio_core_inputs_asyncfifo11_asyncfifo11_readable;
wire [31:0] main_rtio_core_inputs_asyncfifo11_asyncfifo11_din;
wire [31:0] main_rtio_core_inputs_asyncfifo11_asyncfifo11_dout;
wire main_rtio_core_inputs_asyncfifo11_graycounter22_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter22_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo11_graycounter22_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary;
wire main_rtio_core_inputs_asyncfifo11_graycounter23_ce;
(* dont_touch = "true" *) reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter23_q = 3'd0;
wire [2:0] main_rtio_core_inputs_asyncfifo11_graycounter23_q_next;
reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter23_q_binary = 3'd0;
reg [2:0] main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary;
wire [2:0] main_rtio_core_inputs_asyncfifo11_produce_rdomain;
wire [2:0] main_rtio_core_inputs_asyncfifo11_consume_wdomain;
wire [1:0] main_rtio_core_inputs_asyncfifo11_wrport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo11_wrport_dat_r;
wire main_rtio_core_inputs_asyncfifo11_wrport_we;
wire [31:0] main_rtio_core_inputs_asyncfifo11_wrport_dat_w;
wire [1:0] main_rtio_core_inputs_asyncfifo11_rdport_adr;
wire [31:0] main_rtio_core_inputs_asyncfifo11_rdport_dat_r;
wire [31:0] main_rtio_core_inputs_record11_fifo_in_data;
wire [31:0] main_rtio_core_inputs_record11_fifo_out_data;
wire main_rtio_core_inputs_overflow_io11;
wire main_rtio_core_inputs_blindtransfer11_i;
wire main_rtio_core_inputs_blindtransfer11_o;
wire main_rtio_core_inputs_blindtransfer11_ps_i;
wire main_rtio_core_inputs_blindtransfer11_ps_o;
reg main_rtio_core_inputs_blindtransfer11_ps_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer11_ps_toggle_o;
reg main_rtio_core_inputs_blindtransfer11_ps_toggle_o_r = 1'd0;
wire main_rtio_core_inputs_blindtransfer11_ps_ack_i;
wire main_rtio_core_inputs_blindtransfer11_ps_ack_o;
reg main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o;
reg main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_inputs_blindtransfer11_blind = 1'd0;
wire main_rtio_core_inputs_selected11;
reg main_rtio_core_inputs_overflow11 = 1'd0;
wire [1:0] main_rtio_core_inputs_i_status_raw;
reg [63:0] main_rtio_core_inputs_input_timeout = 64'd0;
reg main_rtio_core_inputs_input_pending = 1'd0;
wire main_rtio_core_o_collision_sync_i;
wire main_rtio_core_o_collision_sync_o;
wire [15:0] main_rtio_core_o_collision_sync_data_i;
wire [15:0] main_rtio_core_o_collision_sync_data_o;
wire main_rtio_core_o_collision_sync_ps_i;
wire main_rtio_core_o_collision_sync_ps_o;
reg main_rtio_core_o_collision_sync_ps_toggle_i = 1'd0;
wire main_rtio_core_o_collision_sync_ps_toggle_o;
reg main_rtio_core_o_collision_sync_ps_toggle_o_r = 1'd0;
wire main_rtio_core_o_collision_sync_ps_ack_i;
wire main_rtio_core_o_collision_sync_ps_ack_o;
reg main_rtio_core_o_collision_sync_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_o_collision_sync_ps_ack_toggle_o;
reg main_rtio_core_o_collision_sync_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_o_collision_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_rtio_core_o_collision_sync_bxfer_data = 16'd0;
wire main_rtio_core_o_busy_sync_i;
wire main_rtio_core_o_busy_sync_o;
wire [15:0] main_rtio_core_o_busy_sync_data_i;
wire [15:0] main_rtio_core_o_busy_sync_data_o;
wire main_rtio_core_o_busy_sync_ps_i;
wire main_rtio_core_o_busy_sync_ps_o;
reg main_rtio_core_o_busy_sync_ps_toggle_i = 1'd0;
wire main_rtio_core_o_busy_sync_ps_toggle_o;
reg main_rtio_core_o_busy_sync_ps_toggle_o_r = 1'd0;
wire main_rtio_core_o_busy_sync_ps_ack_i;
wire main_rtio_core_o_busy_sync_ps_ack_o;
reg main_rtio_core_o_busy_sync_ps_ack_toggle_i = 1'd0;
wire main_rtio_core_o_busy_sync_ps_ack_toggle_o;
reg main_rtio_core_o_busy_sync_ps_ack_toggle_o_r = 1'd0;
reg main_rtio_core_o_busy_sync_blind = 1'd0;
(* dont_touch = "true" *) reg [15:0] main_rtio_core_o_busy_sync_bxfer_data = 16'd0;
reg main_rtio_core_o_collision = 1'd0;
reg main_rtio_core_o_busy = 1'd0;
reg main_rtio_core_o_sequence_error = 1'd0;
reg [31:0] main_rtio_target_storage_full = 32'd0;
wire [31:0] main_rtio_target_storage;
reg main_rtio_target_re = 1'd0;
wire main_rtio_now_hi_re;
wire [31:0] main_rtio_now_hi_r;
wire [31:0] main_rtio_now_hi_w;
wire main_rtio_now_lo_re;
wire [31:0] main_rtio_now_lo_r;
wire [31:0] main_rtio_now_lo_w;
reg [511:0] main_rtio_o_data_storage_full = 512'd0;
wire [511:0] main_rtio_o_data_storage;
reg main_rtio_o_data_re = 1'd0;
wire main_rtio_o_data_we;
wire [511:0] main_rtio_o_data_dat_w;
wire [2:0] main_rtio_o_status_status;
reg [63:0] main_rtio_i_timeout_storage_full = 64'd0;
wire [63:0] main_rtio_i_timeout_storage;
reg main_rtio_i_timeout_re = 1'd0;
wire [31:0] main_rtio_i_data_status;
wire [63:0] main_rtio_i_timestamp_status;
wire [3:0] main_rtio_i_status_status;
wire main_rtio_i_overflow_reset_re;
wire main_rtio_i_overflow_reset_r;
reg main_rtio_i_overflow_reset_w = 1'd0;
reg [63:0] main_rtio_counter_status = 64'd0;
wire main_rtio_counter_update_re;
wire main_rtio_counter_update_r;
reg main_rtio_counter_update_w = 1'd0;
reg [1:0] main_rtio_cri_cmd;
wire [23:0] main_rtio_cri_chan_sel;
wire [63:0] main_rtio_cri_o_timestamp;
wire [511:0] main_rtio_cri_o_data;
wire [7:0] main_rtio_cri_o_address;
wire [2:0] main_rtio_cri_o_status;
wire main_rtio_cri_o_buffer_space_valid;
wire [15:0] main_rtio_cri_o_buffer_space;
wire [63:0] main_rtio_cri_i_timeout;
wire [31:0] main_rtio_cri_i_data;
wire [63:0] main_rtio_cri_i_timestamp;
wire [3:0] main_rtio_cri_i_status;
reg [31:0] main_rtio_now_hi_backing = 32'd0;
reg [63:0] main_rtio_now = 64'd0;
wire [29:0] main_interface0_bus_adr;
reg [511:0] main_interface0_bus_dat_w = 512'd0;
wire [511:0] main_interface0_bus_dat_r;
reg [63:0] main_interface0_bus_sel = 64'd0;
wire main_interface0_bus_cyc;
wire main_interface0_bus_stb;
wire main_interface0_bus_ack;
reg main_interface0_bus_we = 1'd0;
reg [2:0] main_interface0_bus_cti = 3'd0;
reg [1:0] main_interface0_bus_bte = 2'd0;
wire main_interface0_bus_err;
wire main_dma_enable_enable_re;
wire main_dma_enable_enable_r;
reg main_dma_enable_enable_w;
reg main_dma_flow_enable;
reg main_dma_dma_sink_stb = 1'd0;
wire main_dma_dma_sink_ack;
reg main_dma_dma_sink_eop = 1'd0;
reg [29:0] main_dma_dma_sink_payload_address = 30'd0;
wire main_dma_dma_source_stb;
wire main_dma_dma_source_ack;
reg main_dma_dma_source_eop = 1'd0;
reg [511:0] main_dma_dma_source_payload_data = 512'd0;
wire main_dma_dma_bus_stb;
reg main_dma_dma_data_reg_loaded = 1'd0;
reg [35:0] main_dma_dma_storage_full = 36'd0;
wire [29:0] main_dma_dma_storage;
reg main_dma_dma_re = 1'd0;
reg main_dma_dma_enable_r = 1'd0;
wire main_dma_rawslicer_sink_stb;
reg main_dma_rawslicer_sink_ack;
wire main_dma_rawslicer_sink_eop;
wire [511:0] main_dma_rawslicer_sink_payload_data;
wire [615:0] main_dma_rawslicer_source;
reg main_dma_rawslicer_source_stb;
reg [6:0] main_dma_rawslicer_source_consume;
reg main_dma_rawslicer_flush;
reg main_dma_rawslicer_flush_done;
reg [1119:0] main_dma_rawslicer_buf = 1120'd0;
reg [7:0] main_dma_rawslicer_level = 8'd0;
reg [7:0] main_dma_rawslicer_next_level;
reg main_dma_rawslicer_load_buf;
reg main_dma_rawslicer_shift_buf;
reg main_dma_reset = 1'd0;
reg main_dma_record_converter_source_stb;
wire main_dma_record_converter_source_ack;
reg main_dma_record_converter_source_eop;
reg [7:0] main_dma_record_converter_source_payload_length = 8'd0;
wire [23:0] main_dma_record_converter_source_payload_channel;
wire [63:0] main_dma_record_converter_source_payload_timestamp;
wire [7:0] main_dma_record_converter_source_payload_address;
reg [511:0] main_dma_record_converter_source_payload_data;
reg main_dma_record_converter_end_marker_found;
reg main_dma_record_converter_flush;
wire [7:0] main_dma_record_converter_record_raw_length;
wire [23:0] main_dma_record_converter_record_raw_channel;
wire [63:0] main_dma_record_converter_record_raw_timestamp;
wire [7:0] main_dma_record_converter_record_raw_address;
wire [511:0] main_dma_record_converter_record_raw_data;
reg [63:0] main_dma_time_offset_storage_full = 64'd0;
wire [63:0] main_dma_time_offset_storage;
reg main_dma_time_offset_re = 1'd0;
reg main_dma_time_offset_source_stb = 1'd0;
wire main_dma_time_offset_source_ack;
reg main_dma_time_offset_source_eop = 1'd0;
reg [7:0] main_dma_time_offset_source_payload_length = 8'd0;
reg [23:0] main_dma_time_offset_source_payload_channel = 24'd0;
reg [63:0] main_dma_time_offset_source_payload_timestamp = 64'd0;
reg [7:0] main_dma_time_offset_source_payload_address = 8'd0;
reg [511:0] main_dma_time_offset_source_payload_data = 512'd0;
wire main_dma_time_offset_sink_stb;
wire main_dma_time_offset_sink_ack;
wire main_dma_time_offset_sink_eop;
wire [7:0] main_dma_time_offset_sink_payload_length;
wire [23:0] main_dma_time_offset_sink_payload_channel;
wire [63:0] main_dma_time_offset_sink_payload_timestamp;
wire [7:0] main_dma_time_offset_sink_payload_address;
wire [511:0] main_dma_time_offset_sink_payload_data;
wire main_dma_cri_master_error_re;
wire [1:0] main_dma_cri_master_error_r;
reg [1:0] main_dma_cri_master_error_w = 2'd0;
reg [23:0] main_dma_cri_master_error_channel_status = 24'd0;
reg [63:0] main_dma_cri_master_error_timestamp_status = 64'd0;
reg [15:0] main_dma_cri_master_error_address_status = 16'd0;
wire main_dma_cri_master_sink_stb;
reg main_dma_cri_master_sink_ack;
wire main_dma_cri_master_sink_eop;
wire [7:0] main_dma_cri_master_sink_payload_length;
wire [23:0] main_dma_cri_master_sink_payload_channel;
wire [63:0] main_dma_cri_master_sink_payload_timestamp;
wire [7:0] main_dma_cri_master_sink_payload_address;
wire [511:0] main_dma_cri_master_sink_payload_data;
reg [1:0] main_dma_cri_master_cri_cmd;
wire [23:0] main_dma_cri_master_cri_chan_sel;
wire [63:0] main_dma_cri_master_cri_o_timestamp;
wire [511:0] main_dma_cri_master_cri_o_data;
wire [7:0] main_dma_cri_master_cri_o_address;
wire [2:0] main_dma_cri_master_cri_o_status;
wire main_dma_cri_master_cri_o_buffer_space_valid;
wire [15:0] main_dma_cri_master_cri_o_buffer_space;
reg [63:0] main_dma_cri_master_cri_i_timeout = 64'd0;
wire [31:0] main_dma_cri_master_cri_i_data;
wire [63:0] main_dma_cri_master_cri_i_timestamp;
wire [3:0] main_dma_cri_master_cri_i_status;
reg main_dma_cri_master_busy;
reg main_dma_cri_master_underflow_trigger;
reg main_dma_cri_master_link_error_trigger;
wire [29:0] main_csrbank0_bus_adr;
wire [31:0] main_csrbank0_bus_dat_w;
reg [31:0] main_csrbank0_bus_dat_r = 32'd0;
wire [3:0] main_csrbank0_bus_sel;
wire main_csrbank0_bus_cyc;
wire main_csrbank0_bus_stb;
reg main_csrbank0_bus_ack = 1'd0;
wire main_csrbank0_bus_we;
wire [2:0] main_csrbank0_bus_cti;
wire [1:0] main_csrbank0_bus_bte;
reg main_csrbank0_bus_err = 1'd0;
wire main_csrbank0_target0_re;
wire [31:0] main_csrbank0_target0_r;
wire [31:0] main_csrbank0_target0_w;
wire main_csrbank0_o_data15_re;
wire [31:0] main_csrbank0_o_data15_r;
wire [31:0] main_csrbank0_o_data15_w;
wire main_csrbank0_o_data14_re;
wire [31:0] main_csrbank0_o_data14_r;
wire [31:0] main_csrbank0_o_data14_w;
wire main_csrbank0_o_data13_re;
wire [31:0] main_csrbank0_o_data13_r;
wire [31:0] main_csrbank0_o_data13_w;
wire main_csrbank0_o_data12_re;
wire [31:0] main_csrbank0_o_data12_r;
wire [31:0] main_csrbank0_o_data12_w;
wire main_csrbank0_o_data11_re;
wire [31:0] main_csrbank0_o_data11_r;
wire [31:0] main_csrbank0_o_data11_w;
wire main_csrbank0_o_data10_re;
wire [31:0] main_csrbank0_o_data10_r;
wire [31:0] main_csrbank0_o_data10_w;
wire main_csrbank0_o_data9_re;
wire [31:0] main_csrbank0_o_data9_r;
wire [31:0] main_csrbank0_o_data9_w;
wire main_csrbank0_o_data8_re;
wire [31:0] main_csrbank0_o_data8_r;
wire [31:0] main_csrbank0_o_data8_w;
wire main_csrbank0_o_data7_re;
wire [31:0] main_csrbank0_o_data7_r;
wire [31:0] main_csrbank0_o_data7_w;
wire main_csrbank0_o_data6_re;
wire [31:0] main_csrbank0_o_data6_r;
wire [31:0] main_csrbank0_o_data6_w;
wire main_csrbank0_o_data5_re;
wire [31:0] main_csrbank0_o_data5_r;
wire [31:0] main_csrbank0_o_data5_w;
wire main_csrbank0_o_data4_re;
wire [31:0] main_csrbank0_o_data4_r;
wire [31:0] main_csrbank0_o_data4_w;
wire main_csrbank0_o_data3_re;
wire [31:0] main_csrbank0_o_data3_r;
wire [31:0] main_csrbank0_o_data3_w;
wire main_csrbank0_o_data2_re;
wire [31:0] main_csrbank0_o_data2_r;
wire [31:0] main_csrbank0_o_data2_w;
wire main_csrbank0_o_data1_re;
wire [31:0] main_csrbank0_o_data1_r;
wire [31:0] main_csrbank0_o_data1_w;
wire main_csrbank0_o_data0_re;
wire [31:0] main_csrbank0_o_data0_r;
wire [31:0] main_csrbank0_o_data0_w;
wire main_csrbank0_o_status_re;
wire [2:0] main_csrbank0_o_status_r;
wire [2:0] main_csrbank0_o_status_w;
wire main_csrbank0_i_timeout1_re;
wire [31:0] main_csrbank0_i_timeout1_r;
wire [31:0] main_csrbank0_i_timeout1_w;
wire main_csrbank0_i_timeout0_re;
wire [31:0] main_csrbank0_i_timeout0_r;
wire [31:0] main_csrbank0_i_timeout0_w;
wire main_csrbank0_i_data_re;
wire [31:0] main_csrbank0_i_data_r;
wire [31:0] main_csrbank0_i_data_w;
wire main_csrbank0_i_timestamp1_re;
wire [31:0] main_csrbank0_i_timestamp1_r;
wire [31:0] main_csrbank0_i_timestamp1_w;
wire main_csrbank0_i_timestamp0_re;
wire [31:0] main_csrbank0_i_timestamp0_r;
wire [31:0] main_csrbank0_i_timestamp0_w;
wire main_csrbank0_i_status_re;
wire [3:0] main_csrbank0_i_status_r;
wire [3:0] main_csrbank0_i_status_w;
wire main_csrbank0_counter1_re;
wire [31:0] main_csrbank0_counter1_r;
wire [31:0] main_csrbank0_counter1_w;
wire main_csrbank0_counter0_re;
wire [31:0] main_csrbank0_counter0_r;
wire [31:0] main_csrbank0_counter0_w;
wire [29:0] main_csrbank1_bus_adr;
wire [31:0] main_csrbank1_bus_dat_w;
reg [31:0] main_csrbank1_bus_dat_r = 32'd0;
wire [3:0] main_csrbank1_bus_sel;
wire main_csrbank1_bus_cyc;
wire main_csrbank1_bus_stb;
reg main_csrbank1_bus_ack = 1'd0;
wire main_csrbank1_bus_we;
wire [2:0] main_csrbank1_bus_cti;
wire [1:0] main_csrbank1_bus_bte;
reg main_csrbank1_bus_err = 1'd0;
wire main_csrbank1_base_address1_re;
wire [3:0] main_csrbank1_base_address1_r;
wire [3:0] main_csrbank1_base_address1_w;
wire main_csrbank1_base_address0_re;
wire [31:0] main_csrbank1_base_address0_r;
wire [31:0] main_csrbank1_base_address0_w;
wire main_csrbank1_time_offset1_re;
wire [31:0] main_csrbank1_time_offset1_r;
wire [31:0] main_csrbank1_time_offset1_w;
wire main_csrbank1_time_offset0_re;
wire [31:0] main_csrbank1_time_offset0_r;
wire [31:0] main_csrbank1_time_offset0_w;
wire main_csrbank1_error_channel_re;
wire [23:0] main_csrbank1_error_channel_r;
wire [23:0] main_csrbank1_error_channel_w;
wire main_csrbank1_error_timestamp1_re;
wire [31:0] main_csrbank1_error_timestamp1_r;
wire [31:0] main_csrbank1_error_timestamp1_w;
wire main_csrbank1_error_timestamp0_re;
wire [31:0] main_csrbank1_error_timestamp0_r;
wire [31:0] main_csrbank1_error_timestamp0_w;
wire main_csrbank1_error_address_re;
wire [15:0] main_csrbank1_error_address_r;
wire [15:0] main_csrbank1_error_address_w;
wire [1:0] main_cri_con_shared_cmd;
wire [23:0] main_cri_con_shared_chan_sel;
wire [63:0] main_cri_con_shared_o_timestamp;
wire [511:0] main_cri_con_shared_o_data;
wire [7:0] main_cri_con_shared_o_address;
reg [2:0] main_cri_con_shared_o_status;
reg main_cri_con_shared_o_buffer_space_valid;
reg [15:0] main_cri_con_shared_o_buffer_space;
wire [63:0] main_cri_con_shared_i_timeout;
reg [31:0] main_cri_con_shared_i_data;
reg [63:0] main_cri_con_shared_i_timestamp;
reg [3:0] main_cri_con_shared_i_status;
reg [1:0] main_cri_con_storage_full = 2'd0;
wire [1:0] main_cri_con_storage;
reg main_cri_con_re = 1'd0;
reg main_cri_con_selected = 1'd0;
wire [29:0] main_csrbank2_bus_adr;
wire [31:0] main_csrbank2_bus_dat_w;
reg [31:0] main_csrbank2_bus_dat_r = 32'd0;
wire [3:0] main_csrbank2_bus_sel;
wire main_csrbank2_bus_cyc;
wire main_csrbank2_bus_stb;
reg main_csrbank2_bus_ack = 1'd0;
wire main_csrbank2_bus_we;
wire [2:0] main_csrbank2_bus_cti;
wire [1:0] main_csrbank2_bus_bte;
reg main_csrbank2_bus_err = 1'd0;
wire main_csrbank2_selected0_re;
wire [1:0] main_csrbank2_selected0_r;
wire [1:0] main_csrbank2_selected0_w;
reg [4:0] main_mon_chan_sel_storage_full = 5'd0;
wire [4:0] main_mon_chan_sel_storage;
reg main_mon_chan_sel_re = 1'd0;
reg [3:0] main_mon_probe_sel_storage_full = 4'd0;
wire [3:0] main_mon_probe_sel_storage;
reg main_mon_probe_sel_re = 1'd0;
wire main_mon_value_update_re;
wire main_mon_value_update_r;
reg main_mon_value_update_w = 1'd0;
reg [31:0] main_mon_status = 32'd0;
wire main_mon_bussynchronizer0_i;
wire main_mon_bussynchronizer0_o;
wire main_mon_bussynchronizer1_i;
wire main_mon_bussynchronizer1_o;
wire main_mon_bussynchronizer2_i;
wire main_mon_bussynchronizer2_o;
wire main_mon_bussynchronizer3_i;
wire main_mon_bussynchronizer3_o;
wire main_mon_bussynchronizer4_i;
wire main_mon_bussynchronizer4_o;
wire main_mon_bussynchronizer5_i;
wire main_mon_bussynchronizer5_o;
wire main_mon_bussynchronizer6_i;
wire main_mon_bussynchronizer6_o;
wire main_mon_bussynchronizer7_i;
wire main_mon_bussynchronizer7_o;
wire main_mon_bussynchronizer8_i;
wire main_mon_bussynchronizer8_o;
wire main_mon_bussynchronizer9_i;
wire main_mon_bussynchronizer9_o;
wire main_mon_bussynchronizer10_i;
wire main_mon_bussynchronizer10_o;
wire main_mon_bussynchronizer11_i;
wire main_mon_bussynchronizer11_o;
wire main_mon_bussynchronizer12_i;
wire main_mon_bussynchronizer12_o;
wire main_mon_bussynchronizer13_i;
wire main_mon_bussynchronizer13_o;
wire main_mon_bussynchronizer14_i;
wire main_mon_bussynchronizer14_o;
wire main_mon_bussynchronizer15_i;
wire main_mon_bussynchronizer15_o;
wire main_mon_bussynchronizer16_i;
wire main_mon_bussynchronizer16_o;
wire main_mon_bussynchronizer17_i;
wire main_mon_bussynchronizer17_o;
wire main_mon_bussynchronizer18_i;
wire main_mon_bussynchronizer18_o;
wire main_mon_bussynchronizer19_i;
wire main_mon_bussynchronizer19_o;
wire main_mon_bussynchronizer20_i;
wire main_mon_bussynchronizer20_o;
wire main_mon_bussynchronizer21_i;
wire main_mon_bussynchronizer21_o;
wire main_mon_bussynchronizer22_i;
wire main_mon_bussynchronizer22_o;
wire main_mon_bussynchronizer23_i;
wire main_mon_bussynchronizer23_o;
wire main_mon_bussynchronizer24_i;
wire main_mon_bussynchronizer24_o;
wire main_mon_bussynchronizer25_i;
wire main_mon_bussynchronizer25_o;
wire main_mon_bussynchronizer26_i;
wire main_mon_bussynchronizer26_o;
wire main_mon_bussynchronizer27_i;
wire main_mon_bussynchronizer27_o;
wire [31:0] main_mon_bussynchronizer28_i;
reg [31:0] main_mon_bussynchronizer28_o = 32'd0;
reg main_mon_bussynchronizer28_starter = 1'd1;
wire main_mon_bussynchronizer28_ping_i;
wire main_mon_bussynchronizer28_ping_o0;
reg main_mon_bussynchronizer28_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer28_ping_toggle_o;
reg main_mon_bussynchronizer28_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer28_ping_o1 = 1'd0;
wire main_mon_bussynchronizer28_pong_i;
wire main_mon_bussynchronizer28_pong_o;
reg main_mon_bussynchronizer28_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer28_pong_toggle_o;
reg main_mon_bussynchronizer28_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer28_wait;
wire main_mon_bussynchronizer28_done;
reg [7:0] main_mon_bussynchronizer28_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer28_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer28_obuffer;
wire [31:0] main_mon_bussynchronizer29_i;
reg [31:0] main_mon_bussynchronizer29_o = 32'd0;
reg main_mon_bussynchronizer29_starter = 1'd1;
wire main_mon_bussynchronizer29_ping_i;
wire main_mon_bussynchronizer29_ping_o0;
reg main_mon_bussynchronizer29_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer29_ping_toggle_o;
reg main_mon_bussynchronizer29_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer29_ping_o1 = 1'd0;
wire main_mon_bussynchronizer29_pong_i;
wire main_mon_bussynchronizer29_pong_o;
reg main_mon_bussynchronizer29_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer29_pong_toggle_o;
reg main_mon_bussynchronizer29_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer29_wait;
wire main_mon_bussynchronizer29_done;
reg [7:0] main_mon_bussynchronizer29_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer29_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer29_obuffer;
wire [31:0] main_mon_bussynchronizer30_i;
reg [31:0] main_mon_bussynchronizer30_o = 32'd0;
reg main_mon_bussynchronizer30_starter = 1'd1;
wire main_mon_bussynchronizer30_ping_i;
wire main_mon_bussynchronizer30_ping_o0;
reg main_mon_bussynchronizer30_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer30_ping_toggle_o;
reg main_mon_bussynchronizer30_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer30_ping_o1 = 1'd0;
wire main_mon_bussynchronizer30_pong_i;
wire main_mon_bussynchronizer30_pong_o;
reg main_mon_bussynchronizer30_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer30_pong_toggle_o;
reg main_mon_bussynchronizer30_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer30_wait;
wire main_mon_bussynchronizer30_done;
reg [7:0] main_mon_bussynchronizer30_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer30_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer30_obuffer;
wire [31:0] main_mon_bussynchronizer31_i;
reg [31:0] main_mon_bussynchronizer31_o = 32'd0;
reg main_mon_bussynchronizer31_starter = 1'd1;
wire main_mon_bussynchronizer31_ping_i;
wire main_mon_bussynchronizer31_ping_o0;
reg main_mon_bussynchronizer31_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer31_ping_toggle_o;
reg main_mon_bussynchronizer31_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer31_ping_o1 = 1'd0;
wire main_mon_bussynchronizer31_pong_i;
wire main_mon_bussynchronizer31_pong_o;
reg main_mon_bussynchronizer31_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer31_pong_toggle_o;
reg main_mon_bussynchronizer31_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer31_wait;
wire main_mon_bussynchronizer31_done;
reg [7:0] main_mon_bussynchronizer31_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer31_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer31_obuffer;
wire [31:0] main_mon_bussynchronizer32_i;
reg [31:0] main_mon_bussynchronizer32_o = 32'd0;
reg main_mon_bussynchronizer32_starter = 1'd1;
wire main_mon_bussynchronizer32_ping_i;
wire main_mon_bussynchronizer32_ping_o0;
reg main_mon_bussynchronizer32_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer32_ping_toggle_o;
reg main_mon_bussynchronizer32_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer32_ping_o1 = 1'd0;
wire main_mon_bussynchronizer32_pong_i;
wire main_mon_bussynchronizer32_pong_o;
reg main_mon_bussynchronizer32_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer32_pong_toggle_o;
reg main_mon_bussynchronizer32_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer32_wait;
wire main_mon_bussynchronizer32_done;
reg [7:0] main_mon_bussynchronizer32_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer32_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer32_obuffer;
wire [31:0] main_mon_bussynchronizer33_i;
reg [31:0] main_mon_bussynchronizer33_o = 32'd0;
reg main_mon_bussynchronizer33_starter = 1'd1;
wire main_mon_bussynchronizer33_ping_i;
wire main_mon_bussynchronizer33_ping_o0;
reg main_mon_bussynchronizer33_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer33_ping_toggle_o;
reg main_mon_bussynchronizer33_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer33_ping_o1 = 1'd0;
wire main_mon_bussynchronizer33_pong_i;
wire main_mon_bussynchronizer33_pong_o;
reg main_mon_bussynchronizer33_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer33_pong_toggle_o;
reg main_mon_bussynchronizer33_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer33_wait;
wire main_mon_bussynchronizer33_done;
reg [7:0] main_mon_bussynchronizer33_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer33_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer33_obuffer;
wire [31:0] main_mon_bussynchronizer34_i;
reg [31:0] main_mon_bussynchronizer34_o = 32'd0;
reg main_mon_bussynchronizer34_starter = 1'd1;
wire main_mon_bussynchronizer34_ping_i;
wire main_mon_bussynchronizer34_ping_o0;
reg main_mon_bussynchronizer34_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer34_ping_toggle_o;
reg main_mon_bussynchronizer34_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer34_ping_o1 = 1'd0;
wire main_mon_bussynchronizer34_pong_i;
wire main_mon_bussynchronizer34_pong_o;
reg main_mon_bussynchronizer34_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer34_pong_toggle_o;
reg main_mon_bussynchronizer34_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer34_wait;
wire main_mon_bussynchronizer34_done;
reg [7:0] main_mon_bussynchronizer34_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer34_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer34_obuffer;
wire [31:0] main_mon_bussynchronizer35_i;
reg [31:0] main_mon_bussynchronizer35_o = 32'd0;
reg main_mon_bussynchronizer35_starter = 1'd1;
wire main_mon_bussynchronizer35_ping_i;
wire main_mon_bussynchronizer35_ping_o0;
reg main_mon_bussynchronizer35_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer35_ping_toggle_o;
reg main_mon_bussynchronizer35_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer35_ping_o1 = 1'd0;
wire main_mon_bussynchronizer35_pong_i;
wire main_mon_bussynchronizer35_pong_o;
reg main_mon_bussynchronizer35_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer35_pong_toggle_o;
reg main_mon_bussynchronizer35_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer35_wait;
wire main_mon_bussynchronizer35_done;
reg [7:0] main_mon_bussynchronizer35_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer35_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer35_obuffer;
wire [31:0] main_mon_bussynchronizer36_i;
reg [31:0] main_mon_bussynchronizer36_o = 32'd0;
reg main_mon_bussynchronizer36_starter = 1'd1;
wire main_mon_bussynchronizer36_ping_i;
wire main_mon_bussynchronizer36_ping_o0;
reg main_mon_bussynchronizer36_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer36_ping_toggle_o;
reg main_mon_bussynchronizer36_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer36_ping_o1 = 1'd0;
wire main_mon_bussynchronizer36_pong_i;
wire main_mon_bussynchronizer36_pong_o;
reg main_mon_bussynchronizer36_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer36_pong_toggle_o;
reg main_mon_bussynchronizer36_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer36_wait;
wire main_mon_bussynchronizer36_done;
reg [7:0] main_mon_bussynchronizer36_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer36_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer36_obuffer;
wire [31:0] main_mon_bussynchronizer37_i;
reg [31:0] main_mon_bussynchronizer37_o = 32'd0;
reg main_mon_bussynchronizer37_starter = 1'd1;
wire main_mon_bussynchronizer37_ping_i;
wire main_mon_bussynchronizer37_ping_o0;
reg main_mon_bussynchronizer37_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer37_ping_toggle_o;
reg main_mon_bussynchronizer37_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer37_ping_o1 = 1'd0;
wire main_mon_bussynchronizer37_pong_i;
wire main_mon_bussynchronizer37_pong_o;
reg main_mon_bussynchronizer37_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer37_pong_toggle_o;
reg main_mon_bussynchronizer37_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer37_wait;
wire main_mon_bussynchronizer37_done;
reg [7:0] main_mon_bussynchronizer37_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer37_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer37_obuffer;
wire [31:0] main_mon_bussynchronizer38_i;
reg [31:0] main_mon_bussynchronizer38_o = 32'd0;
reg main_mon_bussynchronizer38_starter = 1'd1;
wire main_mon_bussynchronizer38_ping_i;
wire main_mon_bussynchronizer38_ping_o0;
reg main_mon_bussynchronizer38_ping_toggle_i = 1'd0;
wire main_mon_bussynchronizer38_ping_toggle_o;
reg main_mon_bussynchronizer38_ping_toggle_o_r = 1'd0;
reg main_mon_bussynchronizer38_ping_o1 = 1'd0;
wire main_mon_bussynchronizer38_pong_i;
wire main_mon_bussynchronizer38_pong_o;
reg main_mon_bussynchronizer38_pong_toggle_i = 1'd0;
wire main_mon_bussynchronizer38_pong_toggle_o;
reg main_mon_bussynchronizer38_pong_toggle_o_r = 1'd0;
wire main_mon_bussynchronizer38_wait;
wire main_mon_bussynchronizer38_done;
reg [7:0] main_mon_bussynchronizer38_count = 8'd128;
(* dont_touch = "true" *) reg [31:0] main_mon_bussynchronizer38_ibuffer = 32'd0;
wire [31:0] main_mon_bussynchronizer38_obuffer;
reg [4:0] main_inj_chan_sel_storage_full = 5'd0;
wire [4:0] main_inj_chan_sel_storage;
reg main_inj_chan_sel_re = 1'd0;
reg [1:0] main_inj_override_sel_storage_full = 2'd0;
wire [1:0] main_inj_override_sel_storage;
reg main_inj_override_sel_re = 1'd0;
wire main_inj_value_re;
wire main_inj_value_r;
wire main_inj_value_w;
reg main_inj_o_sys0 = 1'd0;
reg main_inj_o_sys1 = 1'd0;
reg main_inj_o_sys2 = 1'd0;
reg main_inj_o_sys3 = 1'd0;
reg main_inj_o_sys4 = 1'd0;
reg main_inj_o_sys5 = 1'd0;
reg main_inj_o_sys6 = 1'd0;
reg main_inj_o_sys7 = 1'd0;
reg main_inj_o_sys8 = 1'd0;
reg main_inj_o_sys9 = 1'd0;
reg main_inj_o_sys10 = 1'd0;
reg main_inj_o_sys11 = 1'd0;
reg main_inj_o_sys12 = 1'd0;
reg main_inj_o_sys13 = 1'd0;
reg main_inj_o_sys14 = 1'd0;
reg main_inj_o_sys15 = 1'd0;
reg main_inj_o_sys16 = 1'd0;
reg main_inj_o_sys17 = 1'd0;
reg main_inj_o_sys18 = 1'd0;
reg main_inj_o_sys19 = 1'd0;
reg main_inj_o_sys20 = 1'd0;
reg main_inj_o_sys21 = 1'd0;
reg main_inj_o_sys22 = 1'd0;
reg main_inj_o_sys23 = 1'd0;
reg main_inj_o_sys24 = 1'd0;
reg main_inj_o_sys25 = 1'd0;
reg main_inj_o_sys26 = 1'd0;
reg main_inj_o_sys27 = 1'd0;
reg main_inj_o_sys28 = 1'd0;
reg main_inj_o_sys29 = 1'd0;
reg main_inj_o_sys30 = 1'd0;
reg main_inj_o_sys31 = 1'd0;
reg main_inj_o_sys32 = 1'd0;
reg main_inj_o_sys33 = 1'd0;
reg main_inj_o_sys34 = 1'd0;
reg main_inj_o_sys35 = 1'd0;
reg main_inj_o_sys36 = 1'd0;
reg main_inj_o_sys37 = 1'd0;
reg main_inj_o_sys38 = 1'd0;
reg main_inj_o_sys39 = 1'd0;
reg main_inj_o_sys40 = 1'd0;
reg main_inj_o_sys41 = 1'd0;
reg main_inj_o_sys42 = 1'd0;
reg main_inj_o_sys43 = 1'd0;
reg main_inj_o_sys44 = 1'd0;
reg main_inj_o_sys45 = 1'd0;
reg main_inj_o_sys46 = 1'd0;
reg main_inj_o_sys47 = 1'd0;
reg main_inj_o_sys48 = 1'd0;
reg [29:0] main_interface1_bus_adr = 30'd0;
wire [511:0] main_interface1_bus_dat_w;
wire [511:0] main_interface1_bus_dat_r;
reg [63:0] main_interface1_bus_sel;
wire main_interface1_bus_cyc;
wire main_interface1_bus_stb;
wire main_interface1_bus_ack;
wire main_interface1_bus_we;
reg [2:0] main_interface1_bus_cti = 3'd0;
reg [1:0] main_interface1_bus_bte = 2'd0;
wire main_interface1_bus_err;
reg main_rtio_analyzer_enable_storage_full = 1'd0;
wire main_rtio_analyzer_enable_storage;
reg main_rtio_analyzer_enable_re = 1'd0;
reg main_rtio_analyzer_busy_status = 1'd0;
reg main_rtio_analyzer_message_encoder_source_stb = 1'd0;
wire main_rtio_analyzer_message_encoder_source_ack;
reg main_rtio_analyzer_message_encoder_source_eop = 1'd0;
reg [255:0] main_rtio_analyzer_message_encoder_source_payload_data = 256'd0;
reg main_rtio_analyzer_message_encoder_status = 1'd0;
wire main_rtio_analyzer_message_encoder_overflow_reset_re;
wire main_rtio_analyzer_message_encoder_overflow_reset_r;
reg main_rtio_analyzer_message_encoder_overflow_reset_w = 1'd0;
reg main_rtio_analyzer_message_encoder_read_wait_event_r = 1'd0;
reg main_rtio_analyzer_message_encoder_read_done;
reg main_rtio_analyzer_message_encoder_read_overflow;
wire main_rtio_analyzer_message_encoder_input_output_stb;
reg [1:0] main_rtio_analyzer_message_encoder_input_output_message_type;
wire [29:0] main_rtio_analyzer_message_encoder_input_output_channel;
reg [63:0] main_rtio_analyzer_message_encoder_input_output_timestamp;
wire [63:0] main_rtio_analyzer_message_encoder_input_output_rtio_counter;
wire [31:0] main_rtio_analyzer_message_encoder_input_output_address_padding;
reg [63:0] main_rtio_analyzer_message_encoder_input_output_data;
reg main_rtio_analyzer_message_encoder_exception_stb;
wire [1:0] main_rtio_analyzer_message_encoder_exception_message_type;
wire [29:0] main_rtio_analyzer_message_encoder_exception_channel;
reg [63:0] main_rtio_analyzer_message_encoder_exception_padding0 = 64'd0;
wire [63:0] main_rtio_analyzer_message_encoder_exception_rtio_counter;
reg [7:0] main_rtio_analyzer_message_encoder_exception_exception_type;
reg [87:0] main_rtio_analyzer_message_encoder_exception_padding1 = 88'd0;
reg main_rtio_analyzer_message_encoder_just_written = 1'd0;
wire [1:0] main_rtio_analyzer_message_encoder_stopped_message_type;
reg [93:0] main_rtio_analyzer_message_encoder_stopped_padding0 = 94'd0;
wire [63:0] main_rtio_analyzer_message_encoder_stopped_rtio_counter;
reg [95:0] main_rtio_analyzer_message_encoder_stopped_padding1 = 96'd0;
reg main_rtio_analyzer_message_encoder_enable_r = 1'd0;
reg main_rtio_analyzer_message_encoder_stopping = 1'd0;
wire main_rtio_analyzer_fifo_sink_stb;
wire main_rtio_analyzer_fifo_sink_ack;
wire main_rtio_analyzer_fifo_sink_eop;
wire [255:0] main_rtio_analyzer_fifo_sink_payload_data;
wire main_rtio_analyzer_fifo_source_stb;
wire main_rtio_analyzer_fifo_source_ack;
wire main_rtio_analyzer_fifo_source_eop;
wire [255:0] main_rtio_analyzer_fifo_source_payload_data;
wire main_rtio_analyzer_fifo_re;
reg main_rtio_analyzer_fifo_readable = 1'd0;
wire main_rtio_analyzer_fifo_syncfifo_we;
wire main_rtio_analyzer_fifo_syncfifo_writable;
wire main_rtio_analyzer_fifo_syncfifo_re;
wire main_rtio_analyzer_fifo_syncfifo_readable;
wire [256:0] main_rtio_analyzer_fifo_syncfifo_din;
wire [256:0] main_rtio_analyzer_fifo_syncfifo_dout;
reg [7:0] main_rtio_analyzer_fifo_level0 = 8'd0;
reg main_rtio_analyzer_fifo_replace = 1'd0;
reg [6:0] main_rtio_analyzer_fifo_produce = 7'd0;
reg [6:0] main_rtio_analyzer_fifo_consume = 7'd0;
reg [6:0] main_rtio_analyzer_fifo_wrport_adr;
wire [256:0] main_rtio_analyzer_fifo_wrport_dat_r;
wire main_rtio_analyzer_fifo_wrport_we;
wire [256:0] main_rtio_analyzer_fifo_wrport_dat_w;
wire main_rtio_analyzer_fifo_do_read;
wire [6:0] main_rtio_analyzer_fifo_rdport_adr;
wire [256:0] main_rtio_analyzer_fifo_rdport_dat_r;
wire main_rtio_analyzer_fifo_rdport_re;
wire [7:0] main_rtio_analyzer_fifo_level1;
wire [255:0] main_rtio_analyzer_fifo_fifo_in_payload_data;
wire main_rtio_analyzer_fifo_fifo_in_eop;
wire [255:0] main_rtio_analyzer_fifo_fifo_out_payload_data;
wire main_rtio_analyzer_fifo_fifo_out_eop;
wire main_rtio_analyzer_converter_sink_stb;
wire main_rtio_analyzer_converter_sink_ack;
wire main_rtio_analyzer_converter_sink_eop;
wire [255:0] main_rtio_analyzer_converter_sink_payload_data;
wire main_rtio_analyzer_converter_source_stb;
wire main_rtio_analyzer_converter_source_ack;
reg main_rtio_analyzer_converter_source_eop = 1'd0;
reg [511:0] main_rtio_analyzer_converter_source_payload_data = 512'd0;
reg [1:0] main_rtio_analyzer_converter_source_payload_valid_token_count = 2'd0;
reg main_rtio_analyzer_converter_demux = 1'd0;
wire main_rtio_analyzer_converter_load_part;
reg main_rtio_analyzer_converter_strobe_all = 1'd0;
wire main_rtio_analyzer_dma_reset_re;
wire main_rtio_analyzer_dma_reset_r;
reg main_rtio_analyzer_dma_reset_w = 1'd0;
reg [35:0] main_rtio_analyzer_dma_base_address_storage_full = 36'd0;
wire [29:0] main_rtio_analyzer_dma_base_address_storage;
reg main_rtio_analyzer_dma_base_address_re = 1'd0;
reg [35:0] main_rtio_analyzer_dma_last_address_storage_full = 36'd0;
wire [29:0] main_rtio_analyzer_dma_last_address_storage;
reg main_rtio_analyzer_dma_last_address_re = 1'd0;
wire [63:0] main_rtio_analyzer_dma_status;
wire main_rtio_analyzer_dma_sink_stb;
wire main_rtio_analyzer_dma_sink_ack;
wire main_rtio_analyzer_dma_sink_eop;
wire [511:0] main_rtio_analyzer_dma_sink_payload_data;
wire [1:0] main_rtio_analyzer_dma_sink_payload_valid_token_count;
reg [58:0] main_rtio_analyzer_dma_message_count = 59'd0;
reg main_rtio_analyzer_enable_r = 1'd0;
reg [4:0] builder_minicon_state = 5'd0;
reg [4:0] builder_minicon_next_state;
reg [2:0] builder_fullmemorywe_state = 3'd0;
reg [2:0] builder_fullmemorywe_next_state;
reg [1:0] builder_liteethphygmiimii_state = 2'd0;
reg [1:0] builder_liteethphygmiimii_next_state;
reg builder_liteethmacgap_state = 1'd0;
reg builder_liteethmacgap_next_state;
reg [1:0] builder_liteethmacpreambleinserter_state = 2'd0;
reg [1:0] builder_liteethmacpreambleinserter_next_state;
reg builder_liteethmacpreamblechecker_state = 1'd0;
reg builder_liteethmacpreamblechecker_next_state;
reg [1:0] builder_liteethmaccrc32inserter_state = 2'd0;
reg [1:0] builder_liteethmaccrc32inserter_next_state;
reg [1:0] builder_liteethmaccrc32checker_state = 2'd0;
reg [1:0] builder_liteethmaccrc32checker_next_state;
reg builder_liteethmacpaddinginserter_state = 1'd0;
reg builder_liteethmacpaddinginserter_next_state;
reg [1:0] builder_liteethmacsramwriter_state = 2'd0;
reg [1:0] builder_liteethmacsramwriter_next_state;
reg [31:0] main_writer_errors_status_next_value;
reg main_writer_errors_status_next_value_ce;
reg [1:0] builder_liteethmacsramreader_state = 2'd0;
reg [1:0] builder_liteethmacsramreader_next_state;
wire [29:0] builder_shared_adr;
wire [31:0] builder_shared_dat_w;
wire [31:0] builder_shared_dat_r;
wire [3:0] builder_shared_sel;
wire builder_shared_cyc;
wire builder_shared_stb;
wire builder_shared_ack;
wire builder_shared_we;
wire [2:0] builder_shared_cti;
wire [1:0] builder_shared_bte;
wire builder_shared_err;
wire [1:0] builder_request;
reg builder_grant = 1'd0;
reg [4:0] builder_slave_sel;
reg [4:0] builder_slave_sel_r = 5'd0;
reg [2:0] builder_spimaster0_state = 3'd0;
reg [2:0] builder_spimaster0_next_state;
reg [2:0] builder_spimaster1_state = 3'd0;
reg [2:0] builder_spimaster1_next_state;
reg [2:0] builder_spimaster2_state = 3'd0;
reg [2:0] builder_spimaster2_next_state;
reg [2:0] builder_spimaster3_state = 3'd0;
reg [2:0] builder_spimaster3_next_state;
reg [2:0] builder_spimaster4_state = 3'd0;
reg [2:0] builder_spimaster4_next_state;
reg [2:0] builder_ad9914_state = 3'd0;
reg [2:0] builder_ad9914_next_state;
reg [1:0] builder_resetinserter_state = 2'd0;
reg [1:0] builder_resetinserter_next_state;
reg [1:0] builder_recordconverter_state = 2'd0;
reg [1:0] builder_recordconverter_next_state;
reg [2:0] builder_crimaster_state = 3'd0;
reg [2:0] builder_crimaster_next_state;
reg [2:0] builder_fsm_state = 3'd0;
reg [2:0] builder_fsm_next_state;
wire [1:0] builder_sdram_cpulevel_arbiter_request;
reg builder_sdram_cpulevel_arbiter_grant = 1'd0;
wire [2:0] builder_sdram_native_arbiter_request;
reg [1:0] builder_sdram_native_arbiter_grant = 2'd0;
wire [29:0] builder_nist_clock_shared_adr;
wire [31:0] builder_nist_clock_shared_dat_w;
wire [31:0] builder_nist_clock_shared_dat_r;
wire [3:0] builder_nist_clock_shared_sel;
wire builder_nist_clock_shared_cyc;
wire builder_nist_clock_shared_stb;
wire builder_nist_clock_shared_ack;
wire builder_nist_clock_shared_we;
wire [2:0] builder_nist_clock_shared_cti;
wire [1:0] builder_nist_clock_shared_bte;
wire builder_nist_clock_shared_err;
wire [1:0] builder_nist_clock_request;
reg builder_nist_clock_grant = 1'd0;
reg [5:0] builder_nist_clock_slave_sel;
reg [5:0] builder_nist_clock_slave_sel_r = 6'd0;
wire [13:0] builder_nist_clock_interface0_bank_bus_adr;
wire builder_nist_clock_interface0_bank_bus_we;
wire [7:0] builder_nist_clock_interface0_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface0_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank0_wlevel_en0_re;
wire builder_nist_clock_csrbank0_wlevel_en0_r;
wire builder_nist_clock_csrbank0_wlevel_en0_w;
wire builder_nist_clock_csrbank0_dly_sel0_re;
wire [7:0] builder_nist_clock_csrbank0_dly_sel0_r;
wire [7:0] builder_nist_clock_csrbank0_dly_sel0_w;
wire builder_nist_clock_csrbank0_sel;
wire [13:0] builder_nist_clock_interface1_bank_bus_adr;
wire builder_nist_clock_interface1_bank_bus_we;
wire [7:0] builder_nist_clock_interface1_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface1_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank1_control0_re;
wire [3:0] builder_nist_clock_csrbank1_control0_r;
wire [3:0] builder_nist_clock_csrbank1_control0_w;
wire builder_nist_clock_csrbank1_pi0_command0_re;
wire [5:0] builder_nist_clock_csrbank1_pi0_command0_r;
wire [5:0] builder_nist_clock_csrbank1_pi0_command0_w;
wire builder_nist_clock_csrbank1_pi0_address1_re;
wire [5:0] builder_nist_clock_csrbank1_pi0_address1_r;
wire [5:0] builder_nist_clock_csrbank1_pi0_address1_w;
wire builder_nist_clock_csrbank1_pi0_address0_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_address0_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_address0_w;
wire builder_nist_clock_csrbank1_pi0_baddress0_re;
wire [2:0] builder_nist_clock_csrbank1_pi0_baddress0_r;
wire [2:0] builder_nist_clock_csrbank1_pi0_baddress0_w;
wire builder_nist_clock_csrbank1_pi0_wrdata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata15_w;
wire builder_nist_clock_csrbank1_pi0_wrdata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata14_w;
wire builder_nist_clock_csrbank1_pi0_wrdata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata13_w;
wire builder_nist_clock_csrbank1_pi0_wrdata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata12_w;
wire builder_nist_clock_csrbank1_pi0_wrdata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata11_w;
wire builder_nist_clock_csrbank1_pi0_wrdata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata10_w;
wire builder_nist_clock_csrbank1_pi0_wrdata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata9_w;
wire builder_nist_clock_csrbank1_pi0_wrdata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata8_w;
wire builder_nist_clock_csrbank1_pi0_wrdata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata7_w;
wire builder_nist_clock_csrbank1_pi0_wrdata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata6_w;
wire builder_nist_clock_csrbank1_pi0_wrdata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata5_w;
wire builder_nist_clock_csrbank1_pi0_wrdata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata4_w;
wire builder_nist_clock_csrbank1_pi0_wrdata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata3_w;
wire builder_nist_clock_csrbank1_pi0_wrdata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata2_w;
wire builder_nist_clock_csrbank1_pi0_wrdata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata1_w;
wire builder_nist_clock_csrbank1_pi0_wrdata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_wrdata0_w;
wire builder_nist_clock_csrbank1_pi0_rddata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata15_w;
wire builder_nist_clock_csrbank1_pi0_rddata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata14_w;
wire builder_nist_clock_csrbank1_pi0_rddata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata13_w;
wire builder_nist_clock_csrbank1_pi0_rddata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata12_w;
wire builder_nist_clock_csrbank1_pi0_rddata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata11_w;
wire builder_nist_clock_csrbank1_pi0_rddata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata10_w;
wire builder_nist_clock_csrbank1_pi0_rddata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata9_w;
wire builder_nist_clock_csrbank1_pi0_rddata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata8_w;
wire builder_nist_clock_csrbank1_pi0_rddata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata7_w;
wire builder_nist_clock_csrbank1_pi0_rddata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata6_w;
wire builder_nist_clock_csrbank1_pi0_rddata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata5_w;
wire builder_nist_clock_csrbank1_pi0_rddata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata4_w;
wire builder_nist_clock_csrbank1_pi0_rddata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata3_w;
wire builder_nist_clock_csrbank1_pi0_rddata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata2_w;
wire builder_nist_clock_csrbank1_pi0_rddata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata1_w;
wire builder_nist_clock_csrbank1_pi0_rddata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi0_rddata0_w;
wire builder_nist_clock_csrbank1_pi1_command0_re;
wire [5:0] builder_nist_clock_csrbank1_pi1_command0_r;
wire [5:0] builder_nist_clock_csrbank1_pi1_command0_w;
wire builder_nist_clock_csrbank1_pi1_address1_re;
wire [5:0] builder_nist_clock_csrbank1_pi1_address1_r;
wire [5:0] builder_nist_clock_csrbank1_pi1_address1_w;
wire builder_nist_clock_csrbank1_pi1_address0_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_address0_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_address0_w;
wire builder_nist_clock_csrbank1_pi1_baddress0_re;
wire [2:0] builder_nist_clock_csrbank1_pi1_baddress0_r;
wire [2:0] builder_nist_clock_csrbank1_pi1_baddress0_w;
wire builder_nist_clock_csrbank1_pi1_wrdata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata15_w;
wire builder_nist_clock_csrbank1_pi1_wrdata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata14_w;
wire builder_nist_clock_csrbank1_pi1_wrdata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata13_w;
wire builder_nist_clock_csrbank1_pi1_wrdata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata12_w;
wire builder_nist_clock_csrbank1_pi1_wrdata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata11_w;
wire builder_nist_clock_csrbank1_pi1_wrdata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata10_w;
wire builder_nist_clock_csrbank1_pi1_wrdata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata9_w;
wire builder_nist_clock_csrbank1_pi1_wrdata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata8_w;
wire builder_nist_clock_csrbank1_pi1_wrdata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata7_w;
wire builder_nist_clock_csrbank1_pi1_wrdata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata6_w;
wire builder_nist_clock_csrbank1_pi1_wrdata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata5_w;
wire builder_nist_clock_csrbank1_pi1_wrdata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata4_w;
wire builder_nist_clock_csrbank1_pi1_wrdata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata3_w;
wire builder_nist_clock_csrbank1_pi1_wrdata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata2_w;
wire builder_nist_clock_csrbank1_pi1_wrdata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata1_w;
wire builder_nist_clock_csrbank1_pi1_wrdata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_wrdata0_w;
wire builder_nist_clock_csrbank1_pi1_rddata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata15_w;
wire builder_nist_clock_csrbank1_pi1_rddata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata14_w;
wire builder_nist_clock_csrbank1_pi1_rddata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata13_w;
wire builder_nist_clock_csrbank1_pi1_rddata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata12_w;
wire builder_nist_clock_csrbank1_pi1_rddata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata11_w;
wire builder_nist_clock_csrbank1_pi1_rddata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata10_w;
wire builder_nist_clock_csrbank1_pi1_rddata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata9_w;
wire builder_nist_clock_csrbank1_pi1_rddata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata8_w;
wire builder_nist_clock_csrbank1_pi1_rddata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata7_w;
wire builder_nist_clock_csrbank1_pi1_rddata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata6_w;
wire builder_nist_clock_csrbank1_pi1_rddata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata5_w;
wire builder_nist_clock_csrbank1_pi1_rddata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata4_w;
wire builder_nist_clock_csrbank1_pi1_rddata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata3_w;
wire builder_nist_clock_csrbank1_pi1_rddata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata2_w;
wire builder_nist_clock_csrbank1_pi1_rddata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata1_w;
wire builder_nist_clock_csrbank1_pi1_rddata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi1_rddata0_w;
wire builder_nist_clock_csrbank1_pi2_command0_re;
wire [5:0] builder_nist_clock_csrbank1_pi2_command0_r;
wire [5:0] builder_nist_clock_csrbank1_pi2_command0_w;
wire builder_nist_clock_csrbank1_pi2_address1_re;
wire [5:0] builder_nist_clock_csrbank1_pi2_address1_r;
wire [5:0] builder_nist_clock_csrbank1_pi2_address1_w;
wire builder_nist_clock_csrbank1_pi2_address0_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_address0_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_address0_w;
wire builder_nist_clock_csrbank1_pi2_baddress0_re;
wire [2:0] builder_nist_clock_csrbank1_pi2_baddress0_r;
wire [2:0] builder_nist_clock_csrbank1_pi2_baddress0_w;
wire builder_nist_clock_csrbank1_pi2_wrdata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata15_w;
wire builder_nist_clock_csrbank1_pi2_wrdata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata14_w;
wire builder_nist_clock_csrbank1_pi2_wrdata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata13_w;
wire builder_nist_clock_csrbank1_pi2_wrdata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata12_w;
wire builder_nist_clock_csrbank1_pi2_wrdata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata11_w;
wire builder_nist_clock_csrbank1_pi2_wrdata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata10_w;
wire builder_nist_clock_csrbank1_pi2_wrdata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata9_w;
wire builder_nist_clock_csrbank1_pi2_wrdata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata8_w;
wire builder_nist_clock_csrbank1_pi2_wrdata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata7_w;
wire builder_nist_clock_csrbank1_pi2_wrdata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata6_w;
wire builder_nist_clock_csrbank1_pi2_wrdata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata5_w;
wire builder_nist_clock_csrbank1_pi2_wrdata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata4_w;
wire builder_nist_clock_csrbank1_pi2_wrdata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata3_w;
wire builder_nist_clock_csrbank1_pi2_wrdata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata2_w;
wire builder_nist_clock_csrbank1_pi2_wrdata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata1_w;
wire builder_nist_clock_csrbank1_pi2_wrdata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_wrdata0_w;
wire builder_nist_clock_csrbank1_pi2_rddata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata15_w;
wire builder_nist_clock_csrbank1_pi2_rddata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata14_w;
wire builder_nist_clock_csrbank1_pi2_rddata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata13_w;
wire builder_nist_clock_csrbank1_pi2_rddata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata12_w;
wire builder_nist_clock_csrbank1_pi2_rddata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata11_w;
wire builder_nist_clock_csrbank1_pi2_rddata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata10_w;
wire builder_nist_clock_csrbank1_pi2_rddata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata9_w;
wire builder_nist_clock_csrbank1_pi2_rddata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata8_w;
wire builder_nist_clock_csrbank1_pi2_rddata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata7_w;
wire builder_nist_clock_csrbank1_pi2_rddata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata6_w;
wire builder_nist_clock_csrbank1_pi2_rddata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata5_w;
wire builder_nist_clock_csrbank1_pi2_rddata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata4_w;
wire builder_nist_clock_csrbank1_pi2_rddata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata3_w;
wire builder_nist_clock_csrbank1_pi2_rddata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata2_w;
wire builder_nist_clock_csrbank1_pi2_rddata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata1_w;
wire builder_nist_clock_csrbank1_pi2_rddata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi2_rddata0_w;
wire builder_nist_clock_csrbank1_pi3_command0_re;
wire [5:0] builder_nist_clock_csrbank1_pi3_command0_r;
wire [5:0] builder_nist_clock_csrbank1_pi3_command0_w;
wire builder_nist_clock_csrbank1_pi3_address1_re;
wire [5:0] builder_nist_clock_csrbank1_pi3_address1_r;
wire [5:0] builder_nist_clock_csrbank1_pi3_address1_w;
wire builder_nist_clock_csrbank1_pi3_address0_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_address0_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_address0_w;
wire builder_nist_clock_csrbank1_pi3_baddress0_re;
wire [2:0] builder_nist_clock_csrbank1_pi3_baddress0_r;
wire [2:0] builder_nist_clock_csrbank1_pi3_baddress0_w;
wire builder_nist_clock_csrbank1_pi3_wrdata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata15_w;
wire builder_nist_clock_csrbank1_pi3_wrdata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata14_w;
wire builder_nist_clock_csrbank1_pi3_wrdata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata13_w;
wire builder_nist_clock_csrbank1_pi3_wrdata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata12_w;
wire builder_nist_clock_csrbank1_pi3_wrdata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata11_w;
wire builder_nist_clock_csrbank1_pi3_wrdata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata10_w;
wire builder_nist_clock_csrbank1_pi3_wrdata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata9_w;
wire builder_nist_clock_csrbank1_pi3_wrdata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata8_w;
wire builder_nist_clock_csrbank1_pi3_wrdata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata7_w;
wire builder_nist_clock_csrbank1_pi3_wrdata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata6_w;
wire builder_nist_clock_csrbank1_pi3_wrdata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata5_w;
wire builder_nist_clock_csrbank1_pi3_wrdata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata4_w;
wire builder_nist_clock_csrbank1_pi3_wrdata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata3_w;
wire builder_nist_clock_csrbank1_pi3_wrdata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata2_w;
wire builder_nist_clock_csrbank1_pi3_wrdata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata1_w;
wire builder_nist_clock_csrbank1_pi3_wrdata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_wrdata0_w;
wire builder_nist_clock_csrbank1_pi3_rddata15_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata15_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata15_w;
wire builder_nist_clock_csrbank1_pi3_rddata14_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata14_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata14_w;
wire builder_nist_clock_csrbank1_pi3_rddata13_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata13_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata13_w;
wire builder_nist_clock_csrbank1_pi3_rddata12_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata12_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata12_w;
wire builder_nist_clock_csrbank1_pi3_rddata11_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata11_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata11_w;
wire builder_nist_clock_csrbank1_pi3_rddata10_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata10_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata10_w;
wire builder_nist_clock_csrbank1_pi3_rddata9_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata9_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata9_w;
wire builder_nist_clock_csrbank1_pi3_rddata8_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata8_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata8_w;
wire builder_nist_clock_csrbank1_pi3_rddata7_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata7_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata7_w;
wire builder_nist_clock_csrbank1_pi3_rddata6_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata6_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata6_w;
wire builder_nist_clock_csrbank1_pi3_rddata5_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata5_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata5_w;
wire builder_nist_clock_csrbank1_pi3_rddata4_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata4_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata4_w;
wire builder_nist_clock_csrbank1_pi3_rddata3_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata3_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata3_w;
wire builder_nist_clock_csrbank1_pi3_rddata2_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata2_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata2_w;
wire builder_nist_clock_csrbank1_pi3_rddata1_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata1_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata1_w;
wire builder_nist_clock_csrbank1_pi3_rddata0_re;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata0_r;
wire [7:0] builder_nist_clock_csrbank1_pi3_rddata0_w;
wire builder_nist_clock_csrbank1_sel;
wire [13:0] builder_nist_clock_interface2_bank_bus_adr;
wire builder_nist_clock_interface2_bank_bus_we;
wire [7:0] builder_nist_clock_interface2_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface2_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank2_sram_writer_slot_re;
wire [1:0] builder_nist_clock_csrbank2_sram_writer_slot_r;
wire [1:0] builder_nist_clock_csrbank2_sram_writer_slot_w;
wire builder_nist_clock_csrbank2_sram_writer_length3_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length3_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length3_w;
wire builder_nist_clock_csrbank2_sram_writer_length2_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length2_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length2_w;
wire builder_nist_clock_csrbank2_sram_writer_length1_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length1_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length1_w;
wire builder_nist_clock_csrbank2_sram_writer_length0_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length0_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_length0_w;
wire builder_nist_clock_csrbank2_sram_writer_errors3_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors3_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors3_w;
wire builder_nist_clock_csrbank2_sram_writer_errors2_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors2_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors2_w;
wire builder_nist_clock_csrbank2_sram_writer_errors1_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors1_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors1_w;
wire builder_nist_clock_csrbank2_sram_writer_errors0_re;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors0_r;
wire [7:0] builder_nist_clock_csrbank2_sram_writer_errors0_w;
wire builder_nist_clock_csrbank2_sram_writer_ev_enable0_re;
wire builder_nist_clock_csrbank2_sram_writer_ev_enable0_r;
wire builder_nist_clock_csrbank2_sram_writer_ev_enable0_w;
wire builder_nist_clock_csrbank2_sram_reader_ready_re;
wire builder_nist_clock_csrbank2_sram_reader_ready_r;
wire builder_nist_clock_csrbank2_sram_reader_ready_w;
wire builder_nist_clock_csrbank2_sram_reader_slot0_re;
wire [1:0] builder_nist_clock_csrbank2_sram_reader_slot0_r;
wire [1:0] builder_nist_clock_csrbank2_sram_reader_slot0_w;
wire builder_nist_clock_csrbank2_sram_reader_length1_re;
wire [2:0] builder_nist_clock_csrbank2_sram_reader_length1_r;
wire [2:0] builder_nist_clock_csrbank2_sram_reader_length1_w;
wire builder_nist_clock_csrbank2_sram_reader_length0_re;
wire [7:0] builder_nist_clock_csrbank2_sram_reader_length0_r;
wire [7:0] builder_nist_clock_csrbank2_sram_reader_length0_w;
wire builder_nist_clock_csrbank2_sram_reader_ev_enable0_re;
wire builder_nist_clock_csrbank2_sram_reader_ev_enable0_r;
wire builder_nist_clock_csrbank2_sram_reader_ev_enable0_w;
wire builder_nist_clock_csrbank2_preamble_errors3_re;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors3_r;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors3_w;
wire builder_nist_clock_csrbank2_preamble_errors2_re;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors2_r;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors2_w;
wire builder_nist_clock_csrbank2_preamble_errors1_re;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors1_r;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors1_w;
wire builder_nist_clock_csrbank2_preamble_errors0_re;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors0_r;
wire [7:0] builder_nist_clock_csrbank2_preamble_errors0_w;
wire builder_nist_clock_csrbank2_crc_errors3_re;
wire [7:0] builder_nist_clock_csrbank2_crc_errors3_r;
wire [7:0] builder_nist_clock_csrbank2_crc_errors3_w;
wire builder_nist_clock_csrbank2_crc_errors2_re;
wire [7:0] builder_nist_clock_csrbank2_crc_errors2_r;
wire [7:0] builder_nist_clock_csrbank2_crc_errors2_w;
wire builder_nist_clock_csrbank2_crc_errors1_re;
wire [7:0] builder_nist_clock_csrbank2_crc_errors1_r;
wire [7:0] builder_nist_clock_csrbank2_crc_errors1_w;
wire builder_nist_clock_csrbank2_crc_errors0_re;
wire [7:0] builder_nist_clock_csrbank2_crc_errors0_r;
wire [7:0] builder_nist_clock_csrbank2_crc_errors0_w;
wire builder_nist_clock_csrbank2_sel;
wire [13:0] builder_nist_clock_interface3_bank_bus_adr;
wire builder_nist_clock_interface3_bank_bus_we;
wire [7:0] builder_nist_clock_interface3_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface3_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank3_mode_detection_mode_re;
wire builder_nist_clock_csrbank3_mode_detection_mode_r;
wire builder_nist_clock_csrbank3_mode_detection_mode_w;
wire builder_nist_clock_csrbank3_crg_reset0_re;
wire builder_nist_clock_csrbank3_crg_reset0_r;
wire builder_nist_clock_csrbank3_crg_reset0_w;
wire builder_nist_clock_csrbank3_sel;
wire [13:0] builder_nist_clock_interface4_bank_bus_adr;
wire builder_nist_clock_interface4_bank_bus_we;
wire [7:0] builder_nist_clock_interface4_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface4_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank4_in_re;
wire [1:0] builder_nist_clock_csrbank4_in_r;
wire [1:0] builder_nist_clock_csrbank4_in_w;
wire builder_nist_clock_csrbank4_out0_re;
wire [1:0] builder_nist_clock_csrbank4_out0_r;
wire [1:0] builder_nist_clock_csrbank4_out0_w;
wire builder_nist_clock_csrbank4_oe0_re;
wire [1:0] builder_nist_clock_csrbank4_oe0_r;
wire [1:0] builder_nist_clock_csrbank4_oe0_w;
wire builder_nist_clock_csrbank4_sel;
wire [13:0] builder_nist_clock_interface5_bank_bus_adr;
wire builder_nist_clock_interface5_bank_bus_we;
wire [7:0] builder_nist_clock_interface5_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface5_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank5_address0_re;
wire [7:0] builder_nist_clock_csrbank5_address0_r;
wire [7:0] builder_nist_clock_csrbank5_address0_w;
wire builder_nist_clock_csrbank5_data_re;
wire [7:0] builder_nist_clock_csrbank5_data_r;
wire [7:0] builder_nist_clock_csrbank5_data_w;
wire builder_nist_clock_csrbank5_sel;
wire [13:0] builder_nist_clock_interface6_bank_bus_adr;
wire builder_nist_clock_interface6_bank_bus_we;
wire [7:0] builder_nist_clock_interface6_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface6_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank6_reset0_re;
wire builder_nist_clock_csrbank6_reset0_r;
wire builder_nist_clock_csrbank6_reset0_w;
wire builder_nist_clock_csrbank6_sel;
wire [13:0] builder_nist_clock_interface7_bank_bus_adr;
wire builder_nist_clock_interface7_bank_bus_we;
wire [7:0] builder_nist_clock_interface7_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface7_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank7_out0_re;
wire [1:0] builder_nist_clock_csrbank7_out0_r;
wire [1:0] builder_nist_clock_csrbank7_out0_w;
wire builder_nist_clock_csrbank7_sel;
wire [13:0] builder_nist_clock_interface8_bank_bus_adr;
wire builder_nist_clock_interface8_bank_bus_we;
wire [7:0] builder_nist_clock_interface8_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface8_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank8_enable0_re;
wire builder_nist_clock_csrbank8_enable0_r;
wire builder_nist_clock_csrbank8_enable0_w;
wire builder_nist_clock_csrbank8_busy_re;
wire builder_nist_clock_csrbank8_busy_r;
wire builder_nist_clock_csrbank8_busy_w;
wire builder_nist_clock_csrbank8_message_encoder_overflow_re;
wire builder_nist_clock_csrbank8_message_encoder_overflow_r;
wire builder_nist_clock_csrbank8_message_encoder_overflow_w;
wire builder_nist_clock_csrbank8_dma_base_address4_re;
wire [3:0] builder_nist_clock_csrbank8_dma_base_address4_r;
wire [3:0] builder_nist_clock_csrbank8_dma_base_address4_w;
wire builder_nist_clock_csrbank8_dma_base_address3_re;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address3_r;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address3_w;
wire builder_nist_clock_csrbank8_dma_base_address2_re;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address2_r;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address2_w;
wire builder_nist_clock_csrbank8_dma_base_address1_re;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address1_r;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address1_w;
wire builder_nist_clock_csrbank8_dma_base_address0_re;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address0_r;
wire [7:0] builder_nist_clock_csrbank8_dma_base_address0_w;
wire builder_nist_clock_csrbank8_dma_last_address4_re;
wire [3:0] builder_nist_clock_csrbank8_dma_last_address4_r;
wire [3:0] builder_nist_clock_csrbank8_dma_last_address4_w;
wire builder_nist_clock_csrbank8_dma_last_address3_re;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address3_r;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address3_w;
wire builder_nist_clock_csrbank8_dma_last_address2_re;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address2_r;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address2_w;
wire builder_nist_clock_csrbank8_dma_last_address1_re;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address1_r;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address1_w;
wire builder_nist_clock_csrbank8_dma_last_address0_re;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address0_r;
wire [7:0] builder_nist_clock_csrbank8_dma_last_address0_w;
wire builder_nist_clock_csrbank8_dma_byte_count7_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count7_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count7_w;
wire builder_nist_clock_csrbank8_dma_byte_count6_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count6_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count6_w;
wire builder_nist_clock_csrbank8_dma_byte_count5_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count5_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count5_w;
wire builder_nist_clock_csrbank8_dma_byte_count4_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count4_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count4_w;
wire builder_nist_clock_csrbank8_dma_byte_count3_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count3_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count3_w;
wire builder_nist_clock_csrbank8_dma_byte_count2_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count2_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count2_w;
wire builder_nist_clock_csrbank8_dma_byte_count1_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count1_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count1_w;
wire builder_nist_clock_csrbank8_dma_byte_count0_re;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count0_r;
wire [7:0] builder_nist_clock_csrbank8_dma_byte_count0_w;
wire builder_nist_clock_csrbank8_sel;
wire [13:0] builder_nist_clock_interface9_bank_bus_adr;
wire builder_nist_clock_interface9_bank_bus_we;
wire [7:0] builder_nist_clock_interface9_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface9_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank9_collision_channel1_re;
wire [7:0] builder_nist_clock_csrbank9_collision_channel1_r;
wire [7:0] builder_nist_clock_csrbank9_collision_channel1_w;
wire builder_nist_clock_csrbank9_collision_channel0_re;
wire [7:0] builder_nist_clock_csrbank9_collision_channel0_r;
wire [7:0] builder_nist_clock_csrbank9_collision_channel0_w;
wire builder_nist_clock_csrbank9_busy_channel1_re;
wire [7:0] builder_nist_clock_csrbank9_busy_channel1_r;
wire [7:0] builder_nist_clock_csrbank9_busy_channel1_w;
wire builder_nist_clock_csrbank9_busy_channel0_re;
wire [7:0] builder_nist_clock_csrbank9_busy_channel0_r;
wire [7:0] builder_nist_clock_csrbank9_busy_channel0_w;
wire builder_nist_clock_csrbank9_sequence_error_channel1_re;
wire [7:0] builder_nist_clock_csrbank9_sequence_error_channel1_r;
wire [7:0] builder_nist_clock_csrbank9_sequence_error_channel1_w;
wire builder_nist_clock_csrbank9_sequence_error_channel0_re;
wire [7:0] builder_nist_clock_csrbank9_sequence_error_channel0_r;
wire [7:0] builder_nist_clock_csrbank9_sequence_error_channel0_w;
wire builder_nist_clock_csrbank9_sel;
wire [13:0] builder_nist_clock_interface10_bank_bus_adr;
wire builder_nist_clock_interface10_bank_bus_we;
wire [7:0] builder_nist_clock_interface10_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface10_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank10_clock_sel0_re;
wire builder_nist_clock_csrbank10_clock_sel0_r;
wire builder_nist_clock_csrbank10_clock_sel0_w;
wire builder_nist_clock_csrbank10_pll_reset0_re;
wire builder_nist_clock_csrbank10_pll_reset0_r;
wire builder_nist_clock_csrbank10_pll_reset0_w;
wire builder_nist_clock_csrbank10_pll_locked_re;
wire builder_nist_clock_csrbank10_pll_locked_r;
wire builder_nist_clock_csrbank10_pll_locked_w;
wire builder_nist_clock_csrbank10_sel;
wire [13:0] builder_nist_clock_interface11_bank_bus_adr;
wire builder_nist_clock_interface11_bank_bus_we;
wire [7:0] builder_nist_clock_interface11_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface11_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank11_mon_chan_sel0_re;
wire [4:0] builder_nist_clock_csrbank11_mon_chan_sel0_r;
wire [4:0] builder_nist_clock_csrbank11_mon_chan_sel0_w;
wire builder_nist_clock_csrbank11_mon_probe_sel0_re;
wire [3:0] builder_nist_clock_csrbank11_mon_probe_sel0_r;
wire [3:0] builder_nist_clock_csrbank11_mon_probe_sel0_w;
wire builder_nist_clock_csrbank11_mon_value3_re;
wire [7:0] builder_nist_clock_csrbank11_mon_value3_r;
wire [7:0] builder_nist_clock_csrbank11_mon_value3_w;
wire builder_nist_clock_csrbank11_mon_value2_re;
wire [7:0] builder_nist_clock_csrbank11_mon_value2_r;
wire [7:0] builder_nist_clock_csrbank11_mon_value2_w;
wire builder_nist_clock_csrbank11_mon_value1_re;
wire [7:0] builder_nist_clock_csrbank11_mon_value1_r;
wire [7:0] builder_nist_clock_csrbank11_mon_value1_w;
wire builder_nist_clock_csrbank11_mon_value0_re;
wire [7:0] builder_nist_clock_csrbank11_mon_value0_r;
wire [7:0] builder_nist_clock_csrbank11_mon_value0_w;
wire builder_nist_clock_csrbank11_inj_chan_sel0_re;
wire [4:0] builder_nist_clock_csrbank11_inj_chan_sel0_r;
wire [4:0] builder_nist_clock_csrbank11_inj_chan_sel0_w;
wire builder_nist_clock_csrbank11_inj_override_sel0_re;
wire [1:0] builder_nist_clock_csrbank11_inj_override_sel0_r;
wire [1:0] builder_nist_clock_csrbank11_inj_override_sel0_w;
wire builder_nist_clock_csrbank11_sel;
wire [13:0] builder_nist_clock_interface12_bank_bus_adr;
wire builder_nist_clock_interface12_bank_bus_we;
wire [7:0] builder_nist_clock_interface12_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface12_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank12_bitbang0_re;
wire [3:0] builder_nist_clock_csrbank12_bitbang0_r;
wire [3:0] builder_nist_clock_csrbank12_bitbang0_w;
wire builder_nist_clock_csrbank12_miso_re;
wire builder_nist_clock_csrbank12_miso_r;
wire builder_nist_clock_csrbank12_miso_w;
wire builder_nist_clock_csrbank12_bitbang_en0_re;
wire builder_nist_clock_csrbank12_bitbang_en0_r;
wire builder_nist_clock_csrbank12_bitbang_en0_w;
wire builder_nist_clock_csrbank12_sel;
wire [13:0] builder_nist_clock_interface13_bank_bus_adr;
wire builder_nist_clock_interface13_bank_bus_we;
wire [7:0] builder_nist_clock_interface13_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface13_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank13_load7_re;
wire [7:0] builder_nist_clock_csrbank13_load7_r;
wire [7:0] builder_nist_clock_csrbank13_load7_w;
wire builder_nist_clock_csrbank13_load6_re;
wire [7:0] builder_nist_clock_csrbank13_load6_r;
wire [7:0] builder_nist_clock_csrbank13_load6_w;
wire builder_nist_clock_csrbank13_load5_re;
wire [7:0] builder_nist_clock_csrbank13_load5_r;
wire [7:0] builder_nist_clock_csrbank13_load5_w;
wire builder_nist_clock_csrbank13_load4_re;
wire [7:0] builder_nist_clock_csrbank13_load4_r;
wire [7:0] builder_nist_clock_csrbank13_load4_w;
wire builder_nist_clock_csrbank13_load3_re;
wire [7:0] builder_nist_clock_csrbank13_load3_r;
wire [7:0] builder_nist_clock_csrbank13_load3_w;
wire builder_nist_clock_csrbank13_load2_re;
wire [7:0] builder_nist_clock_csrbank13_load2_r;
wire [7:0] builder_nist_clock_csrbank13_load2_w;
wire builder_nist_clock_csrbank13_load1_re;
wire [7:0] builder_nist_clock_csrbank13_load1_r;
wire [7:0] builder_nist_clock_csrbank13_load1_w;
wire builder_nist_clock_csrbank13_load0_re;
wire [7:0] builder_nist_clock_csrbank13_load0_r;
wire [7:0] builder_nist_clock_csrbank13_load0_w;
wire builder_nist_clock_csrbank13_reload7_re;
wire [7:0] builder_nist_clock_csrbank13_reload7_r;
wire [7:0] builder_nist_clock_csrbank13_reload7_w;
wire builder_nist_clock_csrbank13_reload6_re;
wire [7:0] builder_nist_clock_csrbank13_reload6_r;
wire [7:0] builder_nist_clock_csrbank13_reload6_w;
wire builder_nist_clock_csrbank13_reload5_re;
wire [7:0] builder_nist_clock_csrbank13_reload5_r;
wire [7:0] builder_nist_clock_csrbank13_reload5_w;
wire builder_nist_clock_csrbank13_reload4_re;
wire [7:0] builder_nist_clock_csrbank13_reload4_r;
wire [7:0] builder_nist_clock_csrbank13_reload4_w;
wire builder_nist_clock_csrbank13_reload3_re;
wire [7:0] builder_nist_clock_csrbank13_reload3_r;
wire [7:0] builder_nist_clock_csrbank13_reload3_w;
wire builder_nist_clock_csrbank13_reload2_re;
wire [7:0] builder_nist_clock_csrbank13_reload2_r;
wire [7:0] builder_nist_clock_csrbank13_reload2_w;
wire builder_nist_clock_csrbank13_reload1_re;
wire [7:0] builder_nist_clock_csrbank13_reload1_r;
wire [7:0] builder_nist_clock_csrbank13_reload1_w;
wire builder_nist_clock_csrbank13_reload0_re;
wire [7:0] builder_nist_clock_csrbank13_reload0_r;
wire [7:0] builder_nist_clock_csrbank13_reload0_w;
wire builder_nist_clock_csrbank13_en0_re;
wire builder_nist_clock_csrbank13_en0_r;
wire builder_nist_clock_csrbank13_en0_w;
wire builder_nist_clock_csrbank13_value7_re;
wire [7:0] builder_nist_clock_csrbank13_value7_r;
wire [7:0] builder_nist_clock_csrbank13_value7_w;
wire builder_nist_clock_csrbank13_value6_re;
wire [7:0] builder_nist_clock_csrbank13_value6_r;
wire [7:0] builder_nist_clock_csrbank13_value6_w;
wire builder_nist_clock_csrbank13_value5_re;
wire [7:0] builder_nist_clock_csrbank13_value5_r;
wire [7:0] builder_nist_clock_csrbank13_value5_w;
wire builder_nist_clock_csrbank13_value4_re;
wire [7:0] builder_nist_clock_csrbank13_value4_r;
wire [7:0] builder_nist_clock_csrbank13_value4_w;
wire builder_nist_clock_csrbank13_value3_re;
wire [7:0] builder_nist_clock_csrbank13_value3_r;
wire [7:0] builder_nist_clock_csrbank13_value3_w;
wire builder_nist_clock_csrbank13_value2_re;
wire [7:0] builder_nist_clock_csrbank13_value2_r;
wire [7:0] builder_nist_clock_csrbank13_value2_w;
wire builder_nist_clock_csrbank13_value1_re;
wire [7:0] builder_nist_clock_csrbank13_value1_r;
wire [7:0] builder_nist_clock_csrbank13_value1_w;
wire builder_nist_clock_csrbank13_value0_re;
wire [7:0] builder_nist_clock_csrbank13_value0_r;
wire [7:0] builder_nist_clock_csrbank13_value0_w;
wire builder_nist_clock_csrbank13_ev_enable0_re;
wire builder_nist_clock_csrbank13_ev_enable0_r;
wire builder_nist_clock_csrbank13_ev_enable0_w;
wire builder_nist_clock_csrbank13_sel;
wire [13:0] builder_nist_clock_interface14_bank_bus_adr;
wire builder_nist_clock_interface14_bank_bus_we;
wire [7:0] builder_nist_clock_interface14_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface14_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank14_load7_re;
wire [7:0] builder_nist_clock_csrbank14_load7_r;
wire [7:0] builder_nist_clock_csrbank14_load7_w;
wire builder_nist_clock_csrbank14_load6_re;
wire [7:0] builder_nist_clock_csrbank14_load6_r;
wire [7:0] builder_nist_clock_csrbank14_load6_w;
wire builder_nist_clock_csrbank14_load5_re;
wire [7:0] builder_nist_clock_csrbank14_load5_r;
wire [7:0] builder_nist_clock_csrbank14_load5_w;
wire builder_nist_clock_csrbank14_load4_re;
wire [7:0] builder_nist_clock_csrbank14_load4_r;
wire [7:0] builder_nist_clock_csrbank14_load4_w;
wire builder_nist_clock_csrbank14_load3_re;
wire [7:0] builder_nist_clock_csrbank14_load3_r;
wire [7:0] builder_nist_clock_csrbank14_load3_w;
wire builder_nist_clock_csrbank14_load2_re;
wire [7:0] builder_nist_clock_csrbank14_load2_r;
wire [7:0] builder_nist_clock_csrbank14_load2_w;
wire builder_nist_clock_csrbank14_load1_re;
wire [7:0] builder_nist_clock_csrbank14_load1_r;
wire [7:0] builder_nist_clock_csrbank14_load1_w;
wire builder_nist_clock_csrbank14_load0_re;
wire [7:0] builder_nist_clock_csrbank14_load0_r;
wire [7:0] builder_nist_clock_csrbank14_load0_w;
wire builder_nist_clock_csrbank14_reload7_re;
wire [7:0] builder_nist_clock_csrbank14_reload7_r;
wire [7:0] builder_nist_clock_csrbank14_reload7_w;
wire builder_nist_clock_csrbank14_reload6_re;
wire [7:0] builder_nist_clock_csrbank14_reload6_r;
wire [7:0] builder_nist_clock_csrbank14_reload6_w;
wire builder_nist_clock_csrbank14_reload5_re;
wire [7:0] builder_nist_clock_csrbank14_reload5_r;
wire [7:0] builder_nist_clock_csrbank14_reload5_w;
wire builder_nist_clock_csrbank14_reload4_re;
wire [7:0] builder_nist_clock_csrbank14_reload4_r;
wire [7:0] builder_nist_clock_csrbank14_reload4_w;
wire builder_nist_clock_csrbank14_reload3_re;
wire [7:0] builder_nist_clock_csrbank14_reload3_r;
wire [7:0] builder_nist_clock_csrbank14_reload3_w;
wire builder_nist_clock_csrbank14_reload2_re;
wire [7:0] builder_nist_clock_csrbank14_reload2_r;
wire [7:0] builder_nist_clock_csrbank14_reload2_w;
wire builder_nist_clock_csrbank14_reload1_re;
wire [7:0] builder_nist_clock_csrbank14_reload1_r;
wire [7:0] builder_nist_clock_csrbank14_reload1_w;
wire builder_nist_clock_csrbank14_reload0_re;
wire [7:0] builder_nist_clock_csrbank14_reload0_r;
wire [7:0] builder_nist_clock_csrbank14_reload0_w;
wire builder_nist_clock_csrbank14_en0_re;
wire builder_nist_clock_csrbank14_en0_r;
wire builder_nist_clock_csrbank14_en0_w;
wire builder_nist_clock_csrbank14_value7_re;
wire [7:0] builder_nist_clock_csrbank14_value7_r;
wire [7:0] builder_nist_clock_csrbank14_value7_w;
wire builder_nist_clock_csrbank14_value6_re;
wire [7:0] builder_nist_clock_csrbank14_value6_r;
wire [7:0] builder_nist_clock_csrbank14_value6_w;
wire builder_nist_clock_csrbank14_value5_re;
wire [7:0] builder_nist_clock_csrbank14_value5_r;
wire [7:0] builder_nist_clock_csrbank14_value5_w;
wire builder_nist_clock_csrbank14_value4_re;
wire [7:0] builder_nist_clock_csrbank14_value4_r;
wire [7:0] builder_nist_clock_csrbank14_value4_w;
wire builder_nist_clock_csrbank14_value3_re;
wire [7:0] builder_nist_clock_csrbank14_value3_r;
wire [7:0] builder_nist_clock_csrbank14_value3_w;
wire builder_nist_clock_csrbank14_value2_re;
wire [7:0] builder_nist_clock_csrbank14_value2_r;
wire [7:0] builder_nist_clock_csrbank14_value2_w;
wire builder_nist_clock_csrbank14_value1_re;
wire [7:0] builder_nist_clock_csrbank14_value1_r;
wire [7:0] builder_nist_clock_csrbank14_value1_w;
wire builder_nist_clock_csrbank14_value0_re;
wire [7:0] builder_nist_clock_csrbank14_value0_r;
wire [7:0] builder_nist_clock_csrbank14_value0_w;
wire builder_nist_clock_csrbank14_ev_enable0_re;
wire builder_nist_clock_csrbank14_ev_enable0_r;
wire builder_nist_clock_csrbank14_ev_enable0_w;
wire builder_nist_clock_csrbank14_sel;
wire [13:0] builder_nist_clock_interface15_bank_bus_adr;
wire builder_nist_clock_interface15_bank_bus_we;
wire [7:0] builder_nist_clock_interface15_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface15_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank15_enable_null0_re;
wire builder_nist_clock_csrbank15_enable_null0_r;
wire builder_nist_clock_csrbank15_enable_null0_w;
wire builder_nist_clock_csrbank15_enable_prog0_re;
wire builder_nist_clock_csrbank15_enable_prog0_r;
wire builder_nist_clock_csrbank15_enable_prog0_w;
wire builder_nist_clock_csrbank15_prog_address3_re;
wire [5:0] builder_nist_clock_csrbank15_prog_address3_r;
wire [5:0] builder_nist_clock_csrbank15_prog_address3_w;
wire builder_nist_clock_csrbank15_prog_address2_re;
wire [7:0] builder_nist_clock_csrbank15_prog_address2_r;
wire [7:0] builder_nist_clock_csrbank15_prog_address2_w;
wire builder_nist_clock_csrbank15_prog_address1_re;
wire [7:0] builder_nist_clock_csrbank15_prog_address1_r;
wire [7:0] builder_nist_clock_csrbank15_prog_address1_w;
wire builder_nist_clock_csrbank15_prog_address0_re;
wire [7:0] builder_nist_clock_csrbank15_prog_address0_r;
wire [7:0] builder_nist_clock_csrbank15_prog_address0_w;
wire builder_nist_clock_csrbank15_sel;
wire [13:0] builder_nist_clock_interface16_bank_bus_adr;
wire builder_nist_clock_interface16_bank_bus_we;
wire [7:0] builder_nist_clock_interface16_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface16_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank16_txfull_re;
wire builder_nist_clock_csrbank16_txfull_r;
wire builder_nist_clock_csrbank16_txfull_w;
wire builder_nist_clock_csrbank16_rxempty_re;
wire builder_nist_clock_csrbank16_rxempty_r;
wire builder_nist_clock_csrbank16_rxempty_w;
wire builder_nist_clock_csrbank16_ev_enable0_re;
wire [1:0] builder_nist_clock_csrbank16_ev_enable0_r;
wire [1:0] builder_nist_clock_csrbank16_ev_enable0_w;
wire builder_nist_clock_csrbank16_sel;
wire [13:0] builder_nist_clock_interface17_bank_bus_adr;
wire builder_nist_clock_interface17_bank_bus_we;
wire [7:0] builder_nist_clock_interface17_bank_bus_dat_w;
reg [7:0] builder_nist_clock_interface17_bank_bus_dat_r = 8'd0;
wire builder_nist_clock_csrbank17_tuning_word3_re;
wire [7:0] builder_nist_clock_csrbank17_tuning_word3_r;
wire [7:0] builder_nist_clock_csrbank17_tuning_word3_w;
wire builder_nist_clock_csrbank17_tuning_word2_re;
wire [7:0] builder_nist_clock_csrbank17_tuning_word2_r;
wire [7:0] builder_nist_clock_csrbank17_tuning_word2_w;
wire builder_nist_clock_csrbank17_tuning_word1_re;
wire [7:0] builder_nist_clock_csrbank17_tuning_word1_r;
wire [7:0] builder_nist_clock_csrbank17_tuning_word1_w;
wire builder_nist_clock_csrbank17_tuning_word0_re;
wire [7:0] builder_nist_clock_csrbank17_tuning_word0_r;
wire [7:0] builder_nist_clock_csrbank17_tuning_word0_w;
wire builder_nist_clock_csrbank17_sel;
reg [29:0] builder_comb_rhs_array_muxed0;
reg [31:0] builder_comb_rhs_array_muxed1;
reg [3:0] builder_comb_rhs_array_muxed2;
reg builder_comb_rhs_array_muxed3;
reg builder_comb_rhs_array_muxed4;
reg builder_comb_rhs_array_muxed5;
reg [2:0] builder_comb_rhs_array_muxed6;
reg [1:0] builder_comb_rhs_array_muxed7;
wire builder_comb_lhs_array_muxed;
reg builder_comb_rhs_array_muxed8;
reg [1:0] builder_comb_rhs_array_muxed9;
reg [1:0] builder_comb_rhs_array_muxed10;
reg [23:0] builder_comb_rhs_array_muxed11;
reg [63:0] builder_comb_rhs_array_muxed12;
reg [511:0] builder_comb_rhs_array_muxed13;
reg [7:0] builder_comb_rhs_array_muxed14;
reg [63:0] builder_comb_rhs_array_muxed15;
reg builder_comb_rhs_array_muxed16;
reg builder_comb_rhs_array_muxed17;
reg builder_comb_rhs_array_muxed18;
reg builder_comb_rhs_array_muxed19;
reg builder_comb_rhs_array_muxed20;
reg builder_comb_rhs_array_muxed21;
reg builder_comb_rhs_array_muxed22;
reg builder_comb_rhs_array_muxed23;
reg builder_comb_rhs_array_muxed24;
reg builder_comb_rhs_array_muxed25;
reg builder_comb_rhs_array_muxed26;
reg builder_comb_rhs_array_muxed27;
reg builder_comb_rhs_array_muxed28;
reg builder_comb_rhs_array_muxed29;
reg builder_comb_rhs_array_muxed30;
reg builder_comb_rhs_array_muxed31;
reg builder_comb_rhs_array_muxed32;
reg builder_comb_rhs_array_muxed33;
reg builder_comb_rhs_array_muxed34;
reg builder_comb_rhs_array_muxed35;
reg builder_comb_rhs_array_muxed36;
reg builder_comb_rhs_array_muxed37;
reg builder_comb_rhs_array_muxed38;
reg builder_comb_rhs_array_muxed39;
reg builder_comb_rhs_array_muxed40;
reg builder_comb_rhs_array_muxed41;
reg builder_comb_rhs_array_muxed42;
reg builder_comb_rhs_array_muxed43;
reg builder_comb_rhs_array_muxed44;
reg builder_comb_rhs_array_muxed45;
reg [29:0] builder_comb_rhs_array_muxed46;
reg [31:0] builder_comb_rhs_array_muxed47;
reg [3:0] builder_comb_rhs_array_muxed48;
reg builder_comb_rhs_array_muxed49;
reg builder_comb_rhs_array_muxed50;
reg builder_comb_rhs_array_muxed51;
reg [2:0] builder_comb_rhs_array_muxed52;
reg [1:0] builder_comb_rhs_array_muxed53;
reg [29:0] builder_comb_rhs_array_muxed54;
reg [511:0] builder_comb_rhs_array_muxed55;
reg [63:0] builder_comb_rhs_array_muxed56;
reg builder_comb_rhs_array_muxed57;
reg builder_comb_rhs_array_muxed58;
reg builder_comb_rhs_array_muxed59;
reg [2:0] builder_comb_rhs_array_muxed60;
reg [1:0] builder_comb_rhs_array_muxed61;
reg [29:0] builder_comb_rhs_array_muxed62;
reg [31:0] builder_comb_rhs_array_muxed63;
reg [3:0] builder_comb_rhs_array_muxed64;
reg builder_comb_rhs_array_muxed65;
reg builder_comb_rhs_array_muxed66;
reg builder_comb_rhs_array_muxed67;
reg [2:0] builder_comb_rhs_array_muxed68;
reg [1:0] builder_comb_rhs_array_muxed69;
reg builder_sync_basiclowerer_array_muxed0;
reg builder_sync_basiclowerer_array_muxed1;
reg builder_sync_basiclowerer_array_muxed2;
reg builder_sync_basiclowerer_array_muxed3;
reg builder_sync_basiclowerer_array_muxed4;
reg builder_sync_basiclowerer_array_muxed5;
reg builder_sync_basiclowerer_array_muxed6;
reg builder_sync_basiclowerer_array_muxed7;
reg [7:0] builder_sync_f_t_array_muxed0;
reg [6:0] builder_sync_f_f_array_muxed0;
reg [7:0] builder_sync_f_t_array_muxed1;
reg [6:0] builder_sync_f_f_array_muxed1;
reg [7:0] builder_sync_f_t_array_muxed2;
reg [6:0] builder_sync_f_f_array_muxed2;
reg [7:0] builder_sync_f_t_array_muxed3;
reg [6:0] builder_sync_f_f_array_muxed3;
reg [7:0] builder_sync_f_t_array_muxed4;
reg [6:0] builder_sync_f_f_array_muxed4;
reg [7:0] builder_sync_f_t_array_muxed5;
reg [6:0] builder_sync_f_f_array_muxed5;
reg [7:0] builder_sync_f_t_array_muxed6;
reg [6:0] builder_sync_f_f_array_muxed6;
reg [7:0] builder_sync_f_t_array_muxed7;
reg [6:0] builder_sync_f_f_array_muxed7;
reg [7:0] builder_sync_f_t_array_muxed8;
reg [6:0] builder_sync_f_f_array_muxed8;
reg [7:0] builder_sync_f_t_array_muxed9;
reg [6:0] builder_sync_f_f_array_muxed9;
reg [7:0] builder_sync_f_t_array_muxed10;
reg [6:0] builder_sync_f_f_array_muxed10;
reg [7:0] builder_sync_f_t_array_muxed11;
reg [6:0] builder_sync_f_f_array_muxed11;
reg [7:0] builder_sync_f_t_array_muxed12;
reg [6:0] builder_sync_f_f_array_muxed12;
reg [7:0] builder_sync_f_t_array_muxed13;
reg [6:0] builder_sync_f_f_array_muxed13;
reg [7:0] builder_sync_f_t_array_muxed14;
reg [6:0] builder_sync_f_f_array_muxed14;
reg [7:0] builder_sync_f_t_array_muxed15;
reg [6:0] builder_sync_f_f_array_muxed15;
reg [7:0] builder_sync_f_t_array_muxed16;
reg [6:0] builder_sync_f_f_array_muxed16;
reg [7:0] builder_sync_f_t_array_muxed17;
reg [6:0] builder_sync_f_f_array_muxed17;
reg [7:0] builder_sync_f_t_array_muxed18;
reg [6:0] builder_sync_f_f_array_muxed18;
reg [60:0] builder_sync_rhs_array_muxed0;
reg [60:0] builder_sync_rhs_array_muxed1;
reg [60:0] builder_sync_t_lhs_array_muxed = 61'd0;
reg [31:0] builder_sync_t_rhs_array_muxed0;
reg [64:0] builder_sync_t_rhs_array_muxed1;
reg [31:0] builder_sync_rhs_array_muxed2;
reg [31:0] builder_sync_t_t_array_muxed0 = 32'd0;
reg [31:0] builder_sync_rhs_array_muxed3;
reg [31:0] builder_sync_t_t_array_muxed1 = 32'd0;
reg [31:0] builder_sync_t_rhs_array_muxed2;
reg builder_sync_t_rhs_array_muxed3;
reg builder_sync_t_rhs_array_muxed4;
reg builder_sync_t_rhs_array_muxed5;
reg builder_sync_t_rhs_array_muxed6;
reg builder_sync_t_rhs_array_muxed7;
reg builder_sync_t_rhs_array_muxed8;
reg builder_sync_t_rhs_array_muxed9;
reg builder_sync_t_rhs_array_muxed10;
reg builder_sync_t_rhs_array_muxed11;
reg builder_sync_t_rhs_array_muxed12;
reg builder_sync_t_rhs_array_muxed13;
reg builder_sync_t_rhs_array_muxed14;
reg builder_sync_t_rhs_array_muxed15;
reg builder_sync_t_rhs_array_muxed16;
reg builder_sync_t_rhs_array_muxed17;
reg builder_sync_t_rhs_array_muxed18;
reg builder_sync_t_rhs_array_muxed19;
reg builder_sync_t_rhs_array_muxed20;
reg builder_sync_t_rhs_array_muxed21;
reg builder_sync_t_rhs_array_muxed22;
reg builder_sync_t_rhs_array_muxed23;
reg builder_sync_t_rhs_array_muxed24;
reg builder_sync_t_rhs_array_muxed25;
reg builder_sync_t_rhs_array_muxed26;
reg builder_sync_t_rhs_array_muxed27;
reg builder_sync_t_rhs_array_muxed28;
reg builder_sync_t_rhs_array_muxed29;
reg [31:0] builder_sync_t_rhs_array_muxed30;
reg builder_sync_t_rhs_array_muxed31;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl0_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl0;
wire builder_xilinxasyncresetsynchronizerimpl0_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl1;
wire builder_xilinxasyncresetsynchronizerimpl1_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl1_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl2_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl3_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl2_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl3_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl3_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl4_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl4_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl5_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl5_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl6_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl6_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl7_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] builder_xilinxmultiregimpl7_regs1 = 7'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl8_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl9_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl9_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl4;
wire builder_xilinxasyncresetsynchronizerimpl4_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl10_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl10_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [60:0] builder_xilinxmultiregimpl11_regs0 = 61'd0;
(* async_reg = "true", dont_touch = "true" *) reg [60:0] builder_xilinxmultiregimpl11_regs1 = 61'd0;
wire builder_xilinxasyncresetsynchronizerimpl5_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl6_rst_meta;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl12_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl12_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl13_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl13_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl14_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl14_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl15_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl15_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl16_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl16_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl17_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl17_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl18_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl18_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl19_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl19_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl20_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl20_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl21_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl21_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl22_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl22_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl23_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl23_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl24_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl24_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl25_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl25_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl26_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl26_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl27_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl27_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl28_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl28_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl29_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl29_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl30_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl30_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl31_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl31_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl32_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl32_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl33_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl33_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl34_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl34_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl36_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl36_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl37_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl37_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl38_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl38_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl39_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl39_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl40_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl40_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl41_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl41_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl42_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl42_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl43_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl43_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl44_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl44_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl45_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl45_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl46_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl46_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl47_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl47_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl48_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl48_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl49_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl49_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl50_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl50_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl51_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl51_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl52_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl52_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl53_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] builder_xilinxmultiregimpl53_regs1 = 10'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl54_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl54_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl55_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl55_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl56_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl56_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl57_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl57_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl58_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl58_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl59_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl59_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl60_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl60_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl61_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl61_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl62_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl62_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl63_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl63_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl64_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl64_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl65_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl65_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl66_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl66_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl67_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl67_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl68_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl68_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl69_regs0 = 8'd0;
(* async_reg = "true", dont_touch = "true" *) reg [7:0] builder_xilinxmultiregimpl69_regs1 = 8'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl70_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl70_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl71_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl71_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl72_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl72_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl73_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] builder_xilinxmultiregimpl73_regs1 = 3'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl74_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl74_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl75_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl75_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl76_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl76_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl77_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl77_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl78_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl78_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl79_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl79_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl80_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl80_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl81_regs0 = 16'd0;
(* async_reg = "true", dont_touch = "true" *) reg [15:0] builder_xilinxmultiregimpl81_regs1 = 16'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl82_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl82_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl83_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl83_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl84_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl84_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl85_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl85_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl86_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl86_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl87_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl87_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl88_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl88_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl89_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl89_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl90_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl90_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl91_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl91_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl92_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl92_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl93_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl93_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl94_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl94_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl95_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl95_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl96_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl96_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl97_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl97_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl98_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl98_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl99_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl99_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl100_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl100_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl101_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl101_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl102_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl102_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl103_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl103_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl104_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl104_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl105_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl105_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl106_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl106_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl107_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl107_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl108_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl108_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl109_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl109_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl110_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl110_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl111_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl111_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl112_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl112_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl113_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl113_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl114_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl114_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl115_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl115_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl116_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl116_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl117_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl117_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl118_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl118_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl119_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl119_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl120_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl120_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl121_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl121_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl122_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl122_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl123_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl123_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl124_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl124_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl125_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl125_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl126_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl126_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl127_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl127_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl128_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl128_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl129_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl129_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl130_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl130_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl131_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl131_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl132_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl132_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl133_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl133_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl134_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl134_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl135_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl135_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl136_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl136_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl137_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl137_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl138_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl138_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl139_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl139_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl140_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl140_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl141_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl141_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl142_regs0 = 32'd0;
(* async_reg = "true", dont_touch = "true" *) reg [31:0] builder_xilinxmultiregimpl142_regs1 = 32'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl143_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl143_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl144_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl144_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl145_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl145_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl146_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl146_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl147_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl147_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl148_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl148_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl149_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl149_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl150_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl150_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl151_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl151_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl152_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl152_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl153_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl153_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl154_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl154_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl155_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl155_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl156_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl156_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl157_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl157_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl158_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl158_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl159_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl159_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl160_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl160_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl161_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl161_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl162_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl162_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl163_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl163_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl164_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl164_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl165_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl165_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl166_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl166_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl167_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl167_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl168_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl168_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl169_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl169_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl170_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl170_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl171_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl171_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl172_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl172_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl173_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl173_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl174_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl174_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl175_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl175_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl176_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl176_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl177_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl177_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl178_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl178_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl179_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl179_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl180_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl180_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl181_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl181_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl182_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl182_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl183_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl183_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl184_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl184_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl185_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl185_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl186_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl186_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl187_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl187_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl188_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl188_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl189_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl189_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl190_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl190_regs1 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl191_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_xilinxmultiregimpl191_regs1 = 1'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on

assign main_nist_clock_ddrphy_dfi_p0_address = main_nist_clock_nist_clock_master_p0_address;
assign main_nist_clock_ddrphy_dfi_p0_bank = main_nist_clock_nist_clock_master_p0_bank;
assign main_nist_clock_ddrphy_dfi_p0_cas_n = main_nist_clock_nist_clock_master_p0_cas_n;
assign main_nist_clock_ddrphy_dfi_p0_cs_n = main_nist_clock_nist_clock_master_p0_cs_n;
assign main_nist_clock_ddrphy_dfi_p0_ras_n = main_nist_clock_nist_clock_master_p0_ras_n;
assign main_nist_clock_ddrphy_dfi_p0_we_n = main_nist_clock_nist_clock_master_p0_we_n;
assign main_nist_clock_ddrphy_dfi_p0_cke = main_nist_clock_nist_clock_master_p0_cke;
assign main_nist_clock_ddrphy_dfi_p0_odt = main_nist_clock_nist_clock_master_p0_odt;
assign main_nist_clock_ddrphy_dfi_p0_reset_n = main_nist_clock_nist_clock_master_p0_reset_n;
assign main_nist_clock_ddrphy_dfi_p0_wrdata = main_nist_clock_nist_clock_master_p0_wrdata;
assign main_nist_clock_ddrphy_dfi_p0_wrdata_en = main_nist_clock_nist_clock_master_p0_wrdata_en;
assign main_nist_clock_ddrphy_dfi_p0_wrdata_mask = main_nist_clock_nist_clock_master_p0_wrdata_mask;
assign main_nist_clock_ddrphy_dfi_p0_rddata_en = main_nist_clock_nist_clock_master_p0_rddata_en;
assign main_nist_clock_nist_clock_master_p0_rddata = main_nist_clock_ddrphy_dfi_p0_rddata;
assign main_nist_clock_nist_clock_master_p0_rddata_valid = main_nist_clock_ddrphy_dfi_p0_rddata_valid;
assign main_nist_clock_ddrphy_dfi_p1_address = main_nist_clock_nist_clock_master_p1_address;
assign main_nist_clock_ddrphy_dfi_p1_bank = main_nist_clock_nist_clock_master_p1_bank;
assign main_nist_clock_ddrphy_dfi_p1_cas_n = main_nist_clock_nist_clock_master_p1_cas_n;
assign main_nist_clock_ddrphy_dfi_p1_cs_n = main_nist_clock_nist_clock_master_p1_cs_n;
assign main_nist_clock_ddrphy_dfi_p1_ras_n = main_nist_clock_nist_clock_master_p1_ras_n;
assign main_nist_clock_ddrphy_dfi_p1_we_n = main_nist_clock_nist_clock_master_p1_we_n;
assign main_nist_clock_ddrphy_dfi_p1_cke = main_nist_clock_nist_clock_master_p1_cke;
assign main_nist_clock_ddrphy_dfi_p1_odt = main_nist_clock_nist_clock_master_p1_odt;
assign main_nist_clock_ddrphy_dfi_p1_reset_n = main_nist_clock_nist_clock_master_p1_reset_n;
assign main_nist_clock_ddrphy_dfi_p1_wrdata = main_nist_clock_nist_clock_master_p1_wrdata;
assign main_nist_clock_ddrphy_dfi_p1_wrdata_en = main_nist_clock_nist_clock_master_p1_wrdata_en;
assign main_nist_clock_ddrphy_dfi_p1_wrdata_mask = main_nist_clock_nist_clock_master_p1_wrdata_mask;
assign main_nist_clock_ddrphy_dfi_p1_rddata_en = main_nist_clock_nist_clock_master_p1_rddata_en;
assign main_nist_clock_nist_clock_master_p1_rddata = main_nist_clock_ddrphy_dfi_p1_rddata;
assign main_nist_clock_nist_clock_master_p1_rddata_valid = main_nist_clock_ddrphy_dfi_p1_rddata_valid;
assign main_nist_clock_ddrphy_dfi_p2_address = main_nist_clock_nist_clock_master_p2_address;
assign main_nist_clock_ddrphy_dfi_p2_bank = main_nist_clock_nist_clock_master_p2_bank;
assign main_nist_clock_ddrphy_dfi_p2_cas_n = main_nist_clock_nist_clock_master_p2_cas_n;
assign main_nist_clock_ddrphy_dfi_p2_cs_n = main_nist_clock_nist_clock_master_p2_cs_n;
assign main_nist_clock_ddrphy_dfi_p2_ras_n = main_nist_clock_nist_clock_master_p2_ras_n;
assign main_nist_clock_ddrphy_dfi_p2_we_n = main_nist_clock_nist_clock_master_p2_we_n;
assign main_nist_clock_ddrphy_dfi_p2_cke = main_nist_clock_nist_clock_master_p2_cke;
assign main_nist_clock_ddrphy_dfi_p2_odt = main_nist_clock_nist_clock_master_p2_odt;
assign main_nist_clock_ddrphy_dfi_p2_reset_n = main_nist_clock_nist_clock_master_p2_reset_n;
assign main_nist_clock_ddrphy_dfi_p2_wrdata = main_nist_clock_nist_clock_master_p2_wrdata;
assign main_nist_clock_ddrphy_dfi_p2_wrdata_en = main_nist_clock_nist_clock_master_p2_wrdata_en;
assign main_nist_clock_ddrphy_dfi_p2_wrdata_mask = main_nist_clock_nist_clock_master_p2_wrdata_mask;
assign main_nist_clock_ddrphy_dfi_p2_rddata_en = main_nist_clock_nist_clock_master_p2_rddata_en;
assign main_nist_clock_nist_clock_master_p2_rddata = main_nist_clock_ddrphy_dfi_p2_rddata;
assign main_nist_clock_nist_clock_master_p2_rddata_valid = main_nist_clock_ddrphy_dfi_p2_rddata_valid;
assign main_nist_clock_ddrphy_dfi_p3_address = main_nist_clock_nist_clock_master_p3_address;
assign main_nist_clock_ddrphy_dfi_p3_bank = main_nist_clock_nist_clock_master_p3_bank;
assign main_nist_clock_ddrphy_dfi_p3_cas_n = main_nist_clock_nist_clock_master_p3_cas_n;
assign main_nist_clock_ddrphy_dfi_p3_cs_n = main_nist_clock_nist_clock_master_p3_cs_n;
assign main_nist_clock_ddrphy_dfi_p3_ras_n = main_nist_clock_nist_clock_master_p3_ras_n;
assign main_nist_clock_ddrphy_dfi_p3_we_n = main_nist_clock_nist_clock_master_p3_we_n;
assign main_nist_clock_ddrphy_dfi_p3_cke = main_nist_clock_nist_clock_master_p3_cke;
assign main_nist_clock_ddrphy_dfi_p3_odt = main_nist_clock_nist_clock_master_p3_odt;
assign main_nist_clock_ddrphy_dfi_p3_reset_n = main_nist_clock_nist_clock_master_p3_reset_n;
assign main_nist_clock_ddrphy_dfi_p3_wrdata = main_nist_clock_nist_clock_master_p3_wrdata;
assign main_nist_clock_ddrphy_dfi_p3_wrdata_en = main_nist_clock_nist_clock_master_p3_wrdata_en;
assign main_nist_clock_ddrphy_dfi_p3_wrdata_mask = main_nist_clock_nist_clock_master_p3_wrdata_mask;
assign main_nist_clock_ddrphy_dfi_p3_rddata_en = main_nist_clock_nist_clock_master_p3_rddata_en;
assign main_nist_clock_nist_clock_master_p3_rddata = main_nist_clock_ddrphy_dfi_p3_rddata;
assign main_nist_clock_nist_clock_master_p3_rddata_valid = main_nist_clock_ddrphy_dfi_p3_rddata_valid;
assign main_nist_clock_nist_clock_slave_p0_address = main_nist_clock_nist_clock_sdram_controller_dfi_p0_address;
assign main_nist_clock_nist_clock_slave_p0_bank = main_nist_clock_nist_clock_sdram_controller_dfi_p0_bank;
assign main_nist_clock_nist_clock_slave_p0_cas_n = main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n;
assign main_nist_clock_nist_clock_slave_p0_cs_n = main_nist_clock_nist_clock_sdram_controller_dfi_p0_cs_n;
assign main_nist_clock_nist_clock_slave_p0_ras_n = main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n;
assign main_nist_clock_nist_clock_slave_p0_we_n = main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n;
assign main_nist_clock_nist_clock_slave_p0_cke = main_nist_clock_nist_clock_sdram_controller_dfi_p0_cke;
assign main_nist_clock_nist_clock_slave_p0_odt = main_nist_clock_nist_clock_sdram_controller_dfi_p0_odt;
assign main_nist_clock_nist_clock_slave_p0_reset_n = main_nist_clock_nist_clock_sdram_controller_dfi_p0_reset_n;
assign main_nist_clock_nist_clock_slave_p0_wrdata = main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata;
assign main_nist_clock_nist_clock_slave_p0_wrdata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata_en;
assign main_nist_clock_nist_clock_slave_p0_wrdata_mask = main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata_mask;
assign main_nist_clock_nist_clock_slave_p0_rddata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_en;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata = main_nist_clock_nist_clock_slave_p0_rddata;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_valid = main_nist_clock_nist_clock_slave_p0_rddata_valid;
assign main_nist_clock_nist_clock_slave_p1_address = main_nist_clock_nist_clock_sdram_controller_dfi_p1_address;
assign main_nist_clock_nist_clock_slave_p1_bank = main_nist_clock_nist_clock_sdram_controller_dfi_p1_bank;
assign main_nist_clock_nist_clock_slave_p1_cas_n = main_nist_clock_nist_clock_sdram_controller_dfi_p1_cas_n;
assign main_nist_clock_nist_clock_slave_p1_cs_n = main_nist_clock_nist_clock_sdram_controller_dfi_p1_cs_n;
assign main_nist_clock_nist_clock_slave_p1_ras_n = main_nist_clock_nist_clock_sdram_controller_dfi_p1_ras_n;
assign main_nist_clock_nist_clock_slave_p1_we_n = main_nist_clock_nist_clock_sdram_controller_dfi_p1_we_n;
assign main_nist_clock_nist_clock_slave_p1_cke = main_nist_clock_nist_clock_sdram_controller_dfi_p1_cke;
assign main_nist_clock_nist_clock_slave_p1_odt = main_nist_clock_nist_clock_sdram_controller_dfi_p1_odt;
assign main_nist_clock_nist_clock_slave_p1_reset_n = main_nist_clock_nist_clock_sdram_controller_dfi_p1_reset_n;
assign main_nist_clock_nist_clock_slave_p1_wrdata = main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata;
assign main_nist_clock_nist_clock_slave_p1_wrdata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata_en;
assign main_nist_clock_nist_clock_slave_p1_wrdata_mask = main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata_mask;
assign main_nist_clock_nist_clock_slave_p1_rddata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata_en;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata = main_nist_clock_nist_clock_slave_p1_rddata;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata_valid = main_nist_clock_nist_clock_slave_p1_rddata_valid;
assign main_nist_clock_nist_clock_slave_p2_address = main_nist_clock_nist_clock_sdram_controller_dfi_p2_address;
assign main_nist_clock_nist_clock_slave_p2_bank = main_nist_clock_nist_clock_sdram_controller_dfi_p2_bank;
assign main_nist_clock_nist_clock_slave_p2_cas_n = main_nist_clock_nist_clock_sdram_controller_dfi_p2_cas_n;
assign main_nist_clock_nist_clock_slave_p2_cs_n = main_nist_clock_nist_clock_sdram_controller_dfi_p2_cs_n;
assign main_nist_clock_nist_clock_slave_p2_ras_n = main_nist_clock_nist_clock_sdram_controller_dfi_p2_ras_n;
assign main_nist_clock_nist_clock_slave_p2_we_n = main_nist_clock_nist_clock_sdram_controller_dfi_p2_we_n;
assign main_nist_clock_nist_clock_slave_p2_cke = main_nist_clock_nist_clock_sdram_controller_dfi_p2_cke;
assign main_nist_clock_nist_clock_slave_p2_odt = main_nist_clock_nist_clock_sdram_controller_dfi_p2_odt;
assign main_nist_clock_nist_clock_slave_p2_reset_n = main_nist_clock_nist_clock_sdram_controller_dfi_p2_reset_n;
assign main_nist_clock_nist_clock_slave_p2_wrdata = main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata;
assign main_nist_clock_nist_clock_slave_p2_wrdata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_en;
assign main_nist_clock_nist_clock_slave_p2_wrdata_mask = main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_mask;
assign main_nist_clock_nist_clock_slave_p2_rddata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata_en;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata = main_nist_clock_nist_clock_slave_p2_rddata;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata_valid = main_nist_clock_nist_clock_slave_p2_rddata_valid;
assign main_nist_clock_nist_clock_slave_p3_address = main_nist_clock_nist_clock_sdram_controller_dfi_p3_address;
assign main_nist_clock_nist_clock_slave_p3_bank = main_nist_clock_nist_clock_sdram_controller_dfi_p3_bank;
assign main_nist_clock_nist_clock_slave_p3_cas_n = main_nist_clock_nist_clock_sdram_controller_dfi_p3_cas_n;
assign main_nist_clock_nist_clock_slave_p3_cs_n = main_nist_clock_nist_clock_sdram_controller_dfi_p3_cs_n;
assign main_nist_clock_nist_clock_slave_p3_ras_n = main_nist_clock_nist_clock_sdram_controller_dfi_p3_ras_n;
assign main_nist_clock_nist_clock_slave_p3_we_n = main_nist_clock_nist_clock_sdram_controller_dfi_p3_we_n;
assign main_nist_clock_nist_clock_slave_p3_cke = main_nist_clock_nist_clock_sdram_controller_dfi_p3_cke;
assign main_nist_clock_nist_clock_slave_p3_odt = main_nist_clock_nist_clock_sdram_controller_dfi_p3_odt;
assign main_nist_clock_nist_clock_slave_p3_reset_n = main_nist_clock_nist_clock_sdram_controller_dfi_p3_reset_n;
assign main_nist_clock_nist_clock_slave_p3_wrdata = main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata;
assign main_nist_clock_nist_clock_slave_p3_wrdata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata_en;
assign main_nist_clock_nist_clock_slave_p3_wrdata_mask = main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata_mask;
assign main_nist_clock_nist_clock_slave_p3_rddata_en = main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata_en;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata = main_nist_clock_nist_clock_slave_p3_rddata;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata_valid = main_nist_clock_nist_clock_slave_p3_rddata_valid;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_interrupt <= 32'd0;
	main_nist_clock_nist_clock_interrupt[0] <= main_nist_clock_nist_clock_uart_irq;
	main_nist_clock_nist_clock_interrupt[1] <= main_nist_clock_nist_clock_timer0_irq;
	main_nist_clock_nist_clock_interrupt[2] <= main_ev_irq;
	main_nist_clock_nist_clock_interrupt[3] <= main_irq;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_ibus_adr = main_nist_clock_nist_clock_i_adr_o[31:2];
assign main_nist_clock_nist_clock_dbus_adr = main_nist_clock_nist_clock_d_adr_o[31:2];
assign main_nist_clock_nist_clock_tmpu_adr = main_nist_clock_nist_clock_dbus_adr;
assign main_nist_clock_nist_clock_tmpu_dat_w = main_nist_clock_nist_clock_dbus_dat_w;
assign main_nist_clock_nist_clock_dbus_dat_r = main_nist_clock_nist_clock_tmpu_dat_r;
assign main_nist_clock_nist_clock_tmpu_sel = main_nist_clock_nist_clock_dbus_sel;
assign main_nist_clock_nist_clock_tmpu_cyc = main_nist_clock_nist_clock_dbus_cyc;
assign main_nist_clock_nist_clock_tmpu_stb = main_nist_clock_nist_clock_dbus_stb;
assign main_nist_clock_nist_clock_tmpu_we = main_nist_clock_nist_clock_dbus_we;
assign main_nist_clock_nist_clock_tmpu_cti = main_nist_clock_nist_clock_dbus_cti;
assign main_nist_clock_nist_clock_tmpu_bte = main_nist_clock_nist_clock_dbus_bte;

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_dbus_ack <= 1'd0;
	main_nist_clock_nist_clock_dbus_err <= 1'd0;
	if (main_nist_clock_nist_clock_tmpu_error) begin
		main_nist_clock_nist_clock_dbus_ack <= 1'd0;
		main_nist_clock_nist_clock_dbus_err <= (main_nist_clock_nist_clock_tmpu_ack | main_nist_clock_nist_clock_tmpu_err);
	end else begin
		main_nist_clock_nist_clock_dbus_ack <= main_nist_clock_nist_clock_tmpu_ack;
		main_nist_clock_nist_clock_dbus_err <= main_nist_clock_nist_clock_tmpu_err;
	end
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sram_we <= 4'd0;
	main_nist_clock_nist_clock_sram_we[0] <= (((main_nist_clock_nist_clock_sram_bus_cyc & main_nist_clock_nist_clock_sram_bus_stb) & main_nist_clock_nist_clock_sram_bus_we) & main_nist_clock_nist_clock_sram_bus_sel[0]);
	main_nist_clock_nist_clock_sram_we[1] <= (((main_nist_clock_nist_clock_sram_bus_cyc & main_nist_clock_nist_clock_sram_bus_stb) & main_nist_clock_nist_clock_sram_bus_we) & main_nist_clock_nist_clock_sram_bus_sel[1]);
	main_nist_clock_nist_clock_sram_we[2] <= (((main_nist_clock_nist_clock_sram_bus_cyc & main_nist_clock_nist_clock_sram_bus_stb) & main_nist_clock_nist_clock_sram_bus_we) & main_nist_clock_nist_clock_sram_bus_sel[2]);
	main_nist_clock_nist_clock_sram_we[3] <= (((main_nist_clock_nist_clock_sram_bus_cyc & main_nist_clock_nist_clock_sram_bus_stb) & main_nist_clock_nist_clock_sram_bus_we) & main_nist_clock_nist_clock_sram_bus_sel[3]);
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sram_adr = main_nist_clock_nist_clock_sram_bus_adr[10:0];
assign main_nist_clock_nist_clock_sram_bus_dat_r = main_nist_clock_nist_clock_sram_dat_r;
assign main_nist_clock_nist_clock_sram_dat_w = main_nist_clock_nist_clock_sram_bus_dat_w;
assign main_nist_clock_nist_clock_uart_tx_fifo_sink_stb = main_nist_clock_nist_clock_uart_rxtx_re;
assign main_nist_clock_nist_clock_uart_tx_fifo_sink_payload_data = main_nist_clock_nist_clock_uart_rxtx_r;
assign main_nist_clock_nist_clock_uart_txfull_status = (~main_nist_clock_nist_clock_uart_tx_fifo_sink_ack);
assign main_nist_clock_nist_clock_uart_phy_sink_stb = main_nist_clock_nist_clock_uart_tx_fifo_source_stb;
assign main_nist_clock_nist_clock_uart_tx_fifo_source_ack = main_nist_clock_nist_clock_uart_phy_sink_ack;
assign main_nist_clock_nist_clock_uart_phy_sink_eop = main_nist_clock_nist_clock_uart_tx_fifo_source_eop;
assign main_nist_clock_nist_clock_uart_phy_sink_payload_data = main_nist_clock_nist_clock_uart_tx_fifo_source_payload_data;
assign main_nist_clock_nist_clock_uart_tx_trigger = (~main_nist_clock_nist_clock_uart_tx_fifo_sink_ack);
assign main_nist_clock_nist_clock_uart_rx_fifo_sink_stb = main_nist_clock_nist_clock_uart_phy_source_stb;
assign main_nist_clock_nist_clock_uart_phy_source_ack = main_nist_clock_nist_clock_uart_rx_fifo_sink_ack;
assign main_nist_clock_nist_clock_uart_rx_fifo_sink_eop = main_nist_clock_nist_clock_uart_phy_source_eop;
assign main_nist_clock_nist_clock_uart_rx_fifo_sink_payload_data = main_nist_clock_nist_clock_uart_phy_source_payload_data;
assign main_nist_clock_nist_clock_uart_rxempty_status = (~main_nist_clock_nist_clock_uart_rx_fifo_source_stb);
assign main_nist_clock_nist_clock_uart_rxtx_w = main_nist_clock_nist_clock_uart_rx_fifo_source_payload_data;
assign main_nist_clock_nist_clock_uart_rx_fifo_source_ack = main_nist_clock_nist_clock_uart_rx_clear;
assign main_nist_clock_nist_clock_uart_rx_trigger = (~main_nist_clock_nist_clock_uart_rx_fifo_source_stb);

// synthesis translate_off
reg dummy_d_3;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_tx_clear <= 1'd0;
	if ((main_nist_clock_nist_clock_uart_pending_re & main_nist_clock_nist_clock_uart_pending_r[0])) begin
		main_nist_clock_nist_clock_uart_tx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_3 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_4;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_status_w <= 2'd0;
	main_nist_clock_nist_clock_uart_status_w[0] <= main_nist_clock_nist_clock_uart_tx_status;
	main_nist_clock_nist_clock_uart_status_w[1] <= main_nist_clock_nist_clock_uart_rx_status;
// synthesis translate_off
	dummy_d_4 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_5;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_rx_clear <= 1'd0;
	if ((main_nist_clock_nist_clock_uart_pending_re & main_nist_clock_nist_clock_uart_pending_r[1])) begin
		main_nist_clock_nist_clock_uart_rx_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_5 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_6;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_pending_w <= 2'd0;
	main_nist_clock_nist_clock_uart_pending_w[0] <= main_nist_clock_nist_clock_uart_tx_pending;
	main_nist_clock_nist_clock_uart_pending_w[1] <= main_nist_clock_nist_clock_uart_rx_pending;
// synthesis translate_off
	dummy_d_6 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_uart_irq = ((main_nist_clock_nist_clock_uart_pending_w[0] & main_nist_clock_nist_clock_uart_storage[0]) | (main_nist_clock_nist_clock_uart_pending_w[1] & main_nist_clock_nist_clock_uart_storage[1]));
assign main_nist_clock_nist_clock_uart_tx_status = main_nist_clock_nist_clock_uart_tx_trigger;
assign main_nist_clock_nist_clock_uart_rx_status = main_nist_clock_nist_clock_uart_rx_trigger;
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_din = {main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_eop, main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_payload_data};
assign {main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_eop, main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_payload_data} = main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_dout;
assign main_nist_clock_nist_clock_uart_tx_fifo_sink_ack = main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable;
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_we = main_nist_clock_nist_clock_uart_tx_fifo_sink_stb;
assign main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_eop = main_nist_clock_nist_clock_uart_tx_fifo_sink_eop;
assign main_nist_clock_nist_clock_uart_tx_fifo_fifo_in_payload_data = main_nist_clock_nist_clock_uart_tx_fifo_sink_payload_data;
assign main_nist_clock_nist_clock_uart_tx_fifo_source_stb = main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_readable;
assign main_nist_clock_nist_clock_uart_tx_fifo_source_eop = main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_eop;
assign main_nist_clock_nist_clock_uart_tx_fifo_source_payload_data = main_nist_clock_nist_clock_uart_tx_fifo_fifo_out_payload_data;
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_re = main_nist_clock_nist_clock_uart_tx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_7;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr <= 4'd0;
	if (main_nist_clock_nist_clock_uart_tx_fifo_replace) begin
		main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr <= (main_nist_clock_nist_clock_uart_tx_fifo_produce - 1'd1);
	end else begin
		main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr <= main_nist_clock_nist_clock_uart_tx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_7 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_uart_tx_fifo_wrport_dat_w = main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_din;
assign main_nist_clock_nist_clock_uart_tx_fifo_wrport_we = (main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_we & (main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable | main_nist_clock_nist_clock_uart_tx_fifo_replace));
assign main_nist_clock_nist_clock_uart_tx_fifo_do_read = (main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_readable & main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_re);
assign main_nist_clock_nist_clock_uart_tx_fifo_rdport_adr = main_nist_clock_nist_clock_uart_tx_fifo_consume;
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_dout = main_nist_clock_nist_clock_uart_tx_fifo_rdport_dat_r;
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable = (main_nist_clock_nist_clock_uart_tx_fifo_level != 5'd16);
assign main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_readable = (main_nist_clock_nist_clock_uart_tx_fifo_level != 1'd0);
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_din = {main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_eop, main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_payload_data};
assign {main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_eop, main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_payload_data} = main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_dout;
assign main_nist_clock_nist_clock_uart_rx_fifo_sink_ack = main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable;
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_we = main_nist_clock_nist_clock_uart_rx_fifo_sink_stb;
assign main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_eop = main_nist_clock_nist_clock_uart_rx_fifo_sink_eop;
assign main_nist_clock_nist_clock_uart_rx_fifo_fifo_in_payload_data = main_nist_clock_nist_clock_uart_rx_fifo_sink_payload_data;
assign main_nist_clock_nist_clock_uart_rx_fifo_source_stb = main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_readable;
assign main_nist_clock_nist_clock_uart_rx_fifo_source_eop = main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_eop;
assign main_nist_clock_nist_clock_uart_rx_fifo_source_payload_data = main_nist_clock_nist_clock_uart_rx_fifo_fifo_out_payload_data;
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_re = main_nist_clock_nist_clock_uart_rx_fifo_source_ack;

// synthesis translate_off
reg dummy_d_8;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr <= 4'd0;
	if (main_nist_clock_nist_clock_uart_rx_fifo_replace) begin
		main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr <= (main_nist_clock_nist_clock_uart_rx_fifo_produce - 1'd1);
	end else begin
		main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr <= main_nist_clock_nist_clock_uart_rx_fifo_produce;
	end
// synthesis translate_off
	dummy_d_8 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_uart_rx_fifo_wrport_dat_w = main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_din;
assign main_nist_clock_nist_clock_uart_rx_fifo_wrport_we = (main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_we & (main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable | main_nist_clock_nist_clock_uart_rx_fifo_replace));
assign main_nist_clock_nist_clock_uart_rx_fifo_do_read = (main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_readable & main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_re);
assign main_nist_clock_nist_clock_uart_rx_fifo_rdport_adr = main_nist_clock_nist_clock_uart_rx_fifo_consume;
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_dout = main_nist_clock_nist_clock_uart_rx_fifo_rdport_dat_r;
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable = (main_nist_clock_nist_clock_uart_rx_fifo_level != 5'd16);
assign main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_readable = (main_nist_clock_nist_clock_uart_rx_fifo_level != 1'd0);
assign main_nist_clock_nist_clock_timer0_zero_trigger = (main_nist_clock_nist_clock_timer0_value != 1'd0);
assign main_nist_clock_nist_clock_timer0_eventmanager_status_w = main_nist_clock_nist_clock_timer0_zero_status;

// synthesis translate_off
reg dummy_d_9;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_timer0_zero_clear <= 1'd0;
	if ((main_nist_clock_nist_clock_timer0_eventmanager_pending_re & main_nist_clock_nist_clock_timer0_eventmanager_pending_r)) begin
		main_nist_clock_nist_clock_timer0_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_9 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_timer0_eventmanager_pending_w = main_nist_clock_nist_clock_timer0_zero_pending;
assign main_nist_clock_nist_clock_timer0_irq = (main_nist_clock_nist_clock_timer0_eventmanager_pending_w & main_nist_clock_nist_clock_timer0_eventmanager_storage);
assign main_nist_clock_nist_clock_timer0_zero_status = main_nist_clock_nist_clock_timer0_zero_trigger;

// synthesis translate_off
reg dummy_d_10;
// synthesis translate_on
always @(*) begin
	main_nist_clock_ddrphy_dqs_serdes_pattern <= 8'd0;
	if (main_nist_clock_ddrphy_wlevel_en_storage) begin
		if (main_nist_clock_ddrphy_wlevel_strobe_re) begin
			main_nist_clock_ddrphy_dqs_serdes_pattern <= 1'd1;
		end else begin
			main_nist_clock_ddrphy_dqs_serdes_pattern <= 1'd0;
		end
	end else begin
		main_nist_clock_ddrphy_dqs_serdes_pattern <= 7'd85;
	end
// synthesis translate_off
	dummy_d_10 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_ddrphy_oe = ((main_nist_clock_ddrphy_last_wrdata_en[1] | main_nist_clock_ddrphy_last_wrdata_en[2]) | main_nist_clock_ddrphy_last_wrdata_en[3]);

// synthesis translate_off
reg dummy_d_11;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_inti_p0_rddata <= 128'd0;
	main_nist_clock_nist_clock_inti_p0_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_inti_p1_rddata <= 128'd0;
	main_nist_clock_nist_clock_inti_p1_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_inti_p2_rddata <= 128'd0;
	main_nist_clock_nist_clock_inti_p2_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_inti_p3_rddata <= 128'd0;
	main_nist_clock_nist_clock_inti_p3_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_slave_p0_rddata <= 128'd0;
	main_nist_clock_nist_clock_slave_p0_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_slave_p1_rddata <= 128'd0;
	main_nist_clock_nist_clock_slave_p1_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_slave_p2_rddata <= 128'd0;
	main_nist_clock_nist_clock_slave_p2_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_slave_p3_rddata <= 128'd0;
	main_nist_clock_nist_clock_slave_p3_rddata_valid <= 1'd0;
	main_nist_clock_nist_clock_master_p0_address <= 14'd0;
	main_nist_clock_nist_clock_master_p0_bank <= 3'd0;
	main_nist_clock_nist_clock_master_p0_cas_n <= 1'd1;
	main_nist_clock_nist_clock_master_p0_cs_n <= 1'd1;
	main_nist_clock_nist_clock_master_p0_ras_n <= 1'd1;
	main_nist_clock_nist_clock_master_p0_we_n <= 1'd1;
	main_nist_clock_nist_clock_master_p0_cke <= 1'd0;
	main_nist_clock_nist_clock_master_p0_odt <= 1'd0;
	main_nist_clock_nist_clock_master_p0_reset_n <= 1'd0;
	main_nist_clock_nist_clock_master_p0_wrdata <= 128'd0;
	main_nist_clock_nist_clock_master_p0_wrdata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p0_wrdata_mask <= 16'd0;
	main_nist_clock_nist_clock_master_p0_rddata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p1_address <= 14'd0;
	main_nist_clock_nist_clock_master_p1_bank <= 3'd0;
	main_nist_clock_nist_clock_master_p1_cas_n <= 1'd1;
	main_nist_clock_nist_clock_master_p1_cs_n <= 1'd1;
	main_nist_clock_nist_clock_master_p1_ras_n <= 1'd1;
	main_nist_clock_nist_clock_master_p1_we_n <= 1'd1;
	main_nist_clock_nist_clock_master_p1_cke <= 1'd0;
	main_nist_clock_nist_clock_master_p1_odt <= 1'd0;
	main_nist_clock_nist_clock_master_p1_reset_n <= 1'd0;
	main_nist_clock_nist_clock_master_p1_wrdata <= 128'd0;
	main_nist_clock_nist_clock_master_p1_wrdata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p1_wrdata_mask <= 16'd0;
	main_nist_clock_nist_clock_master_p1_rddata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p2_address <= 14'd0;
	main_nist_clock_nist_clock_master_p2_bank <= 3'd0;
	main_nist_clock_nist_clock_master_p2_cas_n <= 1'd1;
	main_nist_clock_nist_clock_master_p2_cs_n <= 1'd1;
	main_nist_clock_nist_clock_master_p2_ras_n <= 1'd1;
	main_nist_clock_nist_clock_master_p2_we_n <= 1'd1;
	main_nist_clock_nist_clock_master_p2_cke <= 1'd0;
	main_nist_clock_nist_clock_master_p2_odt <= 1'd0;
	main_nist_clock_nist_clock_master_p2_reset_n <= 1'd0;
	main_nist_clock_nist_clock_master_p2_wrdata <= 128'd0;
	main_nist_clock_nist_clock_master_p2_wrdata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p2_wrdata_mask <= 16'd0;
	main_nist_clock_nist_clock_master_p2_rddata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p3_address <= 14'd0;
	main_nist_clock_nist_clock_master_p3_bank <= 3'd0;
	main_nist_clock_nist_clock_master_p3_cas_n <= 1'd1;
	main_nist_clock_nist_clock_master_p3_cs_n <= 1'd1;
	main_nist_clock_nist_clock_master_p3_ras_n <= 1'd1;
	main_nist_clock_nist_clock_master_p3_we_n <= 1'd1;
	main_nist_clock_nist_clock_master_p3_cke <= 1'd0;
	main_nist_clock_nist_clock_master_p3_odt <= 1'd0;
	main_nist_clock_nist_clock_master_p3_reset_n <= 1'd0;
	main_nist_clock_nist_clock_master_p3_wrdata <= 128'd0;
	main_nist_clock_nist_clock_master_p3_wrdata_en <= 1'd0;
	main_nist_clock_nist_clock_master_p3_wrdata_mask <= 16'd0;
	main_nist_clock_nist_clock_master_p3_rddata_en <= 1'd0;
	if (main_nist_clock_nist_clock_storage[0]) begin
		main_nist_clock_nist_clock_master_p0_address <= main_nist_clock_nist_clock_slave_p0_address;
		main_nist_clock_nist_clock_master_p0_bank <= main_nist_clock_nist_clock_slave_p0_bank;
		main_nist_clock_nist_clock_master_p0_cas_n <= main_nist_clock_nist_clock_slave_p0_cas_n;
		main_nist_clock_nist_clock_master_p0_cs_n <= main_nist_clock_nist_clock_slave_p0_cs_n;
		main_nist_clock_nist_clock_master_p0_ras_n <= main_nist_clock_nist_clock_slave_p0_ras_n;
		main_nist_clock_nist_clock_master_p0_we_n <= main_nist_clock_nist_clock_slave_p0_we_n;
		main_nist_clock_nist_clock_master_p0_cke <= main_nist_clock_nist_clock_slave_p0_cke;
		main_nist_clock_nist_clock_master_p0_odt <= main_nist_clock_nist_clock_slave_p0_odt;
		main_nist_clock_nist_clock_master_p0_reset_n <= main_nist_clock_nist_clock_slave_p0_reset_n;
		main_nist_clock_nist_clock_master_p0_wrdata <= main_nist_clock_nist_clock_slave_p0_wrdata;
		main_nist_clock_nist_clock_master_p0_wrdata_en <= main_nist_clock_nist_clock_slave_p0_wrdata_en;
		main_nist_clock_nist_clock_master_p0_wrdata_mask <= main_nist_clock_nist_clock_slave_p0_wrdata_mask;
		main_nist_clock_nist_clock_master_p0_rddata_en <= main_nist_clock_nist_clock_slave_p0_rddata_en;
		main_nist_clock_nist_clock_slave_p0_rddata <= main_nist_clock_nist_clock_master_p0_rddata;
		main_nist_clock_nist_clock_slave_p0_rddata_valid <= main_nist_clock_nist_clock_master_p0_rddata_valid;
		main_nist_clock_nist_clock_master_p1_address <= main_nist_clock_nist_clock_slave_p1_address;
		main_nist_clock_nist_clock_master_p1_bank <= main_nist_clock_nist_clock_slave_p1_bank;
		main_nist_clock_nist_clock_master_p1_cas_n <= main_nist_clock_nist_clock_slave_p1_cas_n;
		main_nist_clock_nist_clock_master_p1_cs_n <= main_nist_clock_nist_clock_slave_p1_cs_n;
		main_nist_clock_nist_clock_master_p1_ras_n <= main_nist_clock_nist_clock_slave_p1_ras_n;
		main_nist_clock_nist_clock_master_p1_we_n <= main_nist_clock_nist_clock_slave_p1_we_n;
		main_nist_clock_nist_clock_master_p1_cke <= main_nist_clock_nist_clock_slave_p1_cke;
		main_nist_clock_nist_clock_master_p1_odt <= main_nist_clock_nist_clock_slave_p1_odt;
		main_nist_clock_nist_clock_master_p1_reset_n <= main_nist_clock_nist_clock_slave_p1_reset_n;
		main_nist_clock_nist_clock_master_p1_wrdata <= main_nist_clock_nist_clock_slave_p1_wrdata;
		main_nist_clock_nist_clock_master_p1_wrdata_en <= main_nist_clock_nist_clock_slave_p1_wrdata_en;
		main_nist_clock_nist_clock_master_p1_wrdata_mask <= main_nist_clock_nist_clock_slave_p1_wrdata_mask;
		main_nist_clock_nist_clock_master_p1_rddata_en <= main_nist_clock_nist_clock_slave_p1_rddata_en;
		main_nist_clock_nist_clock_slave_p1_rddata <= main_nist_clock_nist_clock_master_p1_rddata;
		main_nist_clock_nist_clock_slave_p1_rddata_valid <= main_nist_clock_nist_clock_master_p1_rddata_valid;
		main_nist_clock_nist_clock_master_p2_address <= main_nist_clock_nist_clock_slave_p2_address;
		main_nist_clock_nist_clock_master_p2_bank <= main_nist_clock_nist_clock_slave_p2_bank;
		main_nist_clock_nist_clock_master_p2_cas_n <= main_nist_clock_nist_clock_slave_p2_cas_n;
		main_nist_clock_nist_clock_master_p2_cs_n <= main_nist_clock_nist_clock_slave_p2_cs_n;
		main_nist_clock_nist_clock_master_p2_ras_n <= main_nist_clock_nist_clock_slave_p2_ras_n;
		main_nist_clock_nist_clock_master_p2_we_n <= main_nist_clock_nist_clock_slave_p2_we_n;
		main_nist_clock_nist_clock_master_p2_cke <= main_nist_clock_nist_clock_slave_p2_cke;
		main_nist_clock_nist_clock_master_p2_odt <= main_nist_clock_nist_clock_slave_p2_odt;
		main_nist_clock_nist_clock_master_p2_reset_n <= main_nist_clock_nist_clock_slave_p2_reset_n;
		main_nist_clock_nist_clock_master_p2_wrdata <= main_nist_clock_nist_clock_slave_p2_wrdata;
		main_nist_clock_nist_clock_master_p2_wrdata_en <= main_nist_clock_nist_clock_slave_p2_wrdata_en;
		main_nist_clock_nist_clock_master_p2_wrdata_mask <= main_nist_clock_nist_clock_slave_p2_wrdata_mask;
		main_nist_clock_nist_clock_master_p2_rddata_en <= main_nist_clock_nist_clock_slave_p2_rddata_en;
		main_nist_clock_nist_clock_slave_p2_rddata <= main_nist_clock_nist_clock_master_p2_rddata;
		main_nist_clock_nist_clock_slave_p2_rddata_valid <= main_nist_clock_nist_clock_master_p2_rddata_valid;
		main_nist_clock_nist_clock_master_p3_address <= main_nist_clock_nist_clock_slave_p3_address;
		main_nist_clock_nist_clock_master_p3_bank <= main_nist_clock_nist_clock_slave_p3_bank;
		main_nist_clock_nist_clock_master_p3_cas_n <= main_nist_clock_nist_clock_slave_p3_cas_n;
		main_nist_clock_nist_clock_master_p3_cs_n <= main_nist_clock_nist_clock_slave_p3_cs_n;
		main_nist_clock_nist_clock_master_p3_ras_n <= main_nist_clock_nist_clock_slave_p3_ras_n;
		main_nist_clock_nist_clock_master_p3_we_n <= main_nist_clock_nist_clock_slave_p3_we_n;
		main_nist_clock_nist_clock_master_p3_cke <= main_nist_clock_nist_clock_slave_p3_cke;
		main_nist_clock_nist_clock_master_p3_odt <= main_nist_clock_nist_clock_slave_p3_odt;
		main_nist_clock_nist_clock_master_p3_reset_n <= main_nist_clock_nist_clock_slave_p3_reset_n;
		main_nist_clock_nist_clock_master_p3_wrdata <= main_nist_clock_nist_clock_slave_p3_wrdata;
		main_nist_clock_nist_clock_master_p3_wrdata_en <= main_nist_clock_nist_clock_slave_p3_wrdata_en;
		main_nist_clock_nist_clock_master_p3_wrdata_mask <= main_nist_clock_nist_clock_slave_p3_wrdata_mask;
		main_nist_clock_nist_clock_master_p3_rddata_en <= main_nist_clock_nist_clock_slave_p3_rddata_en;
		main_nist_clock_nist_clock_slave_p3_rddata <= main_nist_clock_nist_clock_master_p3_rddata;
		main_nist_clock_nist_clock_slave_p3_rddata_valid <= main_nist_clock_nist_clock_master_p3_rddata_valid;
	end else begin
		main_nist_clock_nist_clock_master_p0_address <= main_nist_clock_nist_clock_inti_p0_address;
		main_nist_clock_nist_clock_master_p0_bank <= main_nist_clock_nist_clock_inti_p0_bank;
		main_nist_clock_nist_clock_master_p0_cas_n <= main_nist_clock_nist_clock_inti_p0_cas_n;
		main_nist_clock_nist_clock_master_p0_cs_n <= main_nist_clock_nist_clock_inti_p0_cs_n;
		main_nist_clock_nist_clock_master_p0_ras_n <= main_nist_clock_nist_clock_inti_p0_ras_n;
		main_nist_clock_nist_clock_master_p0_we_n <= main_nist_clock_nist_clock_inti_p0_we_n;
		main_nist_clock_nist_clock_master_p0_cke <= main_nist_clock_nist_clock_inti_p0_cke;
		main_nist_clock_nist_clock_master_p0_odt <= main_nist_clock_nist_clock_inti_p0_odt;
		main_nist_clock_nist_clock_master_p0_reset_n <= main_nist_clock_nist_clock_inti_p0_reset_n;
		main_nist_clock_nist_clock_master_p0_wrdata <= main_nist_clock_nist_clock_inti_p0_wrdata;
		main_nist_clock_nist_clock_master_p0_wrdata_en <= main_nist_clock_nist_clock_inti_p0_wrdata_en;
		main_nist_clock_nist_clock_master_p0_wrdata_mask <= main_nist_clock_nist_clock_inti_p0_wrdata_mask;
		main_nist_clock_nist_clock_master_p0_rddata_en <= main_nist_clock_nist_clock_inti_p0_rddata_en;
		main_nist_clock_nist_clock_inti_p0_rddata <= main_nist_clock_nist_clock_master_p0_rddata;
		main_nist_clock_nist_clock_inti_p0_rddata_valid <= main_nist_clock_nist_clock_master_p0_rddata_valid;
		main_nist_clock_nist_clock_master_p1_address <= main_nist_clock_nist_clock_inti_p1_address;
		main_nist_clock_nist_clock_master_p1_bank <= main_nist_clock_nist_clock_inti_p1_bank;
		main_nist_clock_nist_clock_master_p1_cas_n <= main_nist_clock_nist_clock_inti_p1_cas_n;
		main_nist_clock_nist_clock_master_p1_cs_n <= main_nist_clock_nist_clock_inti_p1_cs_n;
		main_nist_clock_nist_clock_master_p1_ras_n <= main_nist_clock_nist_clock_inti_p1_ras_n;
		main_nist_clock_nist_clock_master_p1_we_n <= main_nist_clock_nist_clock_inti_p1_we_n;
		main_nist_clock_nist_clock_master_p1_cke <= main_nist_clock_nist_clock_inti_p1_cke;
		main_nist_clock_nist_clock_master_p1_odt <= main_nist_clock_nist_clock_inti_p1_odt;
		main_nist_clock_nist_clock_master_p1_reset_n <= main_nist_clock_nist_clock_inti_p1_reset_n;
		main_nist_clock_nist_clock_master_p1_wrdata <= main_nist_clock_nist_clock_inti_p1_wrdata;
		main_nist_clock_nist_clock_master_p1_wrdata_en <= main_nist_clock_nist_clock_inti_p1_wrdata_en;
		main_nist_clock_nist_clock_master_p1_wrdata_mask <= main_nist_clock_nist_clock_inti_p1_wrdata_mask;
		main_nist_clock_nist_clock_master_p1_rddata_en <= main_nist_clock_nist_clock_inti_p1_rddata_en;
		main_nist_clock_nist_clock_inti_p1_rddata <= main_nist_clock_nist_clock_master_p1_rddata;
		main_nist_clock_nist_clock_inti_p1_rddata_valid <= main_nist_clock_nist_clock_master_p1_rddata_valid;
		main_nist_clock_nist_clock_master_p2_address <= main_nist_clock_nist_clock_inti_p2_address;
		main_nist_clock_nist_clock_master_p2_bank <= main_nist_clock_nist_clock_inti_p2_bank;
		main_nist_clock_nist_clock_master_p2_cas_n <= main_nist_clock_nist_clock_inti_p2_cas_n;
		main_nist_clock_nist_clock_master_p2_cs_n <= main_nist_clock_nist_clock_inti_p2_cs_n;
		main_nist_clock_nist_clock_master_p2_ras_n <= main_nist_clock_nist_clock_inti_p2_ras_n;
		main_nist_clock_nist_clock_master_p2_we_n <= main_nist_clock_nist_clock_inti_p2_we_n;
		main_nist_clock_nist_clock_master_p2_cke <= main_nist_clock_nist_clock_inti_p2_cke;
		main_nist_clock_nist_clock_master_p2_odt <= main_nist_clock_nist_clock_inti_p2_odt;
		main_nist_clock_nist_clock_master_p2_reset_n <= main_nist_clock_nist_clock_inti_p2_reset_n;
		main_nist_clock_nist_clock_master_p2_wrdata <= main_nist_clock_nist_clock_inti_p2_wrdata;
		main_nist_clock_nist_clock_master_p2_wrdata_en <= main_nist_clock_nist_clock_inti_p2_wrdata_en;
		main_nist_clock_nist_clock_master_p2_wrdata_mask <= main_nist_clock_nist_clock_inti_p2_wrdata_mask;
		main_nist_clock_nist_clock_master_p2_rddata_en <= main_nist_clock_nist_clock_inti_p2_rddata_en;
		main_nist_clock_nist_clock_inti_p2_rddata <= main_nist_clock_nist_clock_master_p2_rddata;
		main_nist_clock_nist_clock_inti_p2_rddata_valid <= main_nist_clock_nist_clock_master_p2_rddata_valid;
		main_nist_clock_nist_clock_master_p3_address <= main_nist_clock_nist_clock_inti_p3_address;
		main_nist_clock_nist_clock_master_p3_bank <= main_nist_clock_nist_clock_inti_p3_bank;
		main_nist_clock_nist_clock_master_p3_cas_n <= main_nist_clock_nist_clock_inti_p3_cas_n;
		main_nist_clock_nist_clock_master_p3_cs_n <= main_nist_clock_nist_clock_inti_p3_cs_n;
		main_nist_clock_nist_clock_master_p3_ras_n <= main_nist_clock_nist_clock_inti_p3_ras_n;
		main_nist_clock_nist_clock_master_p3_we_n <= main_nist_clock_nist_clock_inti_p3_we_n;
		main_nist_clock_nist_clock_master_p3_cke <= main_nist_clock_nist_clock_inti_p3_cke;
		main_nist_clock_nist_clock_master_p3_odt <= main_nist_clock_nist_clock_inti_p3_odt;
		main_nist_clock_nist_clock_master_p3_reset_n <= main_nist_clock_nist_clock_inti_p3_reset_n;
		main_nist_clock_nist_clock_master_p3_wrdata <= main_nist_clock_nist_clock_inti_p3_wrdata;
		main_nist_clock_nist_clock_master_p3_wrdata_en <= main_nist_clock_nist_clock_inti_p3_wrdata_en;
		main_nist_clock_nist_clock_master_p3_wrdata_mask <= main_nist_clock_nist_clock_inti_p3_wrdata_mask;
		main_nist_clock_nist_clock_master_p3_rddata_en <= main_nist_clock_nist_clock_inti_p3_rddata_en;
		main_nist_clock_nist_clock_inti_p3_rddata <= main_nist_clock_nist_clock_master_p3_rddata;
		main_nist_clock_nist_clock_inti_p3_rddata_valid <= main_nist_clock_nist_clock_master_p3_rddata_valid;
	end
// synthesis translate_off
	dummy_d_11 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_inti_p0_cke = main_nist_clock_nist_clock_storage[1];
assign main_nist_clock_nist_clock_inti_p1_cke = main_nist_clock_nist_clock_storage[1];
assign main_nist_clock_nist_clock_inti_p2_cke = main_nist_clock_nist_clock_storage[1];
assign main_nist_clock_nist_clock_inti_p3_cke = main_nist_clock_nist_clock_storage[1];
assign main_nist_clock_nist_clock_inti_p0_odt = main_nist_clock_nist_clock_storage[2];
assign main_nist_clock_nist_clock_inti_p1_odt = main_nist_clock_nist_clock_storage[2];
assign main_nist_clock_nist_clock_inti_p2_odt = main_nist_clock_nist_clock_storage[2];
assign main_nist_clock_nist_clock_inti_p3_odt = main_nist_clock_nist_clock_storage[2];
assign main_nist_clock_nist_clock_inti_p0_reset_n = main_nist_clock_nist_clock_storage[3];
assign main_nist_clock_nist_clock_inti_p1_reset_n = main_nist_clock_nist_clock_storage[3];
assign main_nist_clock_nist_clock_inti_p2_reset_n = main_nist_clock_nist_clock_storage[3];
assign main_nist_clock_nist_clock_inti_p3_reset_n = main_nist_clock_nist_clock_storage[3];

// synthesis translate_off
reg dummy_d_12;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_inti_p0_cas_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p0_cs_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p0_ras_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p0_we_n <= 1'd1;
	if (main_nist_clock_nist_clock_phaseinjector0_command_issue_re) begin
		main_nist_clock_nist_clock_inti_p0_cs_n <= (~main_nist_clock_nist_clock_phaseinjector0_command_storage[0]);
		main_nist_clock_nist_clock_inti_p0_we_n <= (~main_nist_clock_nist_clock_phaseinjector0_command_storage[1]);
		main_nist_clock_nist_clock_inti_p0_cas_n <= (~main_nist_clock_nist_clock_phaseinjector0_command_storage[2]);
		main_nist_clock_nist_clock_inti_p0_ras_n <= (~main_nist_clock_nist_clock_phaseinjector0_command_storage[3]);
	end else begin
		main_nist_clock_nist_clock_inti_p0_cs_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p0_we_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p0_cas_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p0_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_12 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_inti_p0_address = main_nist_clock_nist_clock_phaseinjector0_address_storage;
assign main_nist_clock_nist_clock_inti_p0_bank = main_nist_clock_nist_clock_phaseinjector0_baddress_storage;
assign main_nist_clock_nist_clock_inti_p0_wrdata_en = (main_nist_clock_nist_clock_phaseinjector0_command_issue_re & main_nist_clock_nist_clock_phaseinjector0_command_storage[4]);
assign main_nist_clock_nist_clock_inti_p0_rddata_en = (main_nist_clock_nist_clock_phaseinjector0_command_issue_re & main_nist_clock_nist_clock_phaseinjector0_command_storage[5]);
assign main_nist_clock_nist_clock_inti_p0_wrdata = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage;
assign main_nist_clock_nist_clock_inti_p0_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_13;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_inti_p1_cas_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p1_cs_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p1_ras_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p1_we_n <= 1'd1;
	if (main_nist_clock_nist_clock_phaseinjector1_command_issue_re) begin
		main_nist_clock_nist_clock_inti_p1_cs_n <= (~main_nist_clock_nist_clock_phaseinjector1_command_storage[0]);
		main_nist_clock_nist_clock_inti_p1_we_n <= (~main_nist_clock_nist_clock_phaseinjector1_command_storage[1]);
		main_nist_clock_nist_clock_inti_p1_cas_n <= (~main_nist_clock_nist_clock_phaseinjector1_command_storage[2]);
		main_nist_clock_nist_clock_inti_p1_ras_n <= (~main_nist_clock_nist_clock_phaseinjector1_command_storage[3]);
	end else begin
		main_nist_clock_nist_clock_inti_p1_cs_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p1_we_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p1_cas_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p1_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_13 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_inti_p1_address = main_nist_clock_nist_clock_phaseinjector1_address_storage;
assign main_nist_clock_nist_clock_inti_p1_bank = main_nist_clock_nist_clock_phaseinjector1_baddress_storage;
assign main_nist_clock_nist_clock_inti_p1_wrdata_en = (main_nist_clock_nist_clock_phaseinjector1_command_issue_re & main_nist_clock_nist_clock_phaseinjector1_command_storage[4]);
assign main_nist_clock_nist_clock_inti_p1_rddata_en = (main_nist_clock_nist_clock_phaseinjector1_command_issue_re & main_nist_clock_nist_clock_phaseinjector1_command_storage[5]);
assign main_nist_clock_nist_clock_inti_p1_wrdata = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage;
assign main_nist_clock_nist_clock_inti_p1_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_14;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_inti_p2_cas_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p2_cs_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p2_ras_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p2_we_n <= 1'd1;
	if (main_nist_clock_nist_clock_phaseinjector2_command_issue_re) begin
		main_nist_clock_nist_clock_inti_p2_cs_n <= (~main_nist_clock_nist_clock_phaseinjector2_command_storage[0]);
		main_nist_clock_nist_clock_inti_p2_we_n <= (~main_nist_clock_nist_clock_phaseinjector2_command_storage[1]);
		main_nist_clock_nist_clock_inti_p2_cas_n <= (~main_nist_clock_nist_clock_phaseinjector2_command_storage[2]);
		main_nist_clock_nist_clock_inti_p2_ras_n <= (~main_nist_clock_nist_clock_phaseinjector2_command_storage[3]);
	end else begin
		main_nist_clock_nist_clock_inti_p2_cs_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p2_we_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p2_cas_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p2_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_14 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_inti_p2_address = main_nist_clock_nist_clock_phaseinjector2_address_storage;
assign main_nist_clock_nist_clock_inti_p2_bank = main_nist_clock_nist_clock_phaseinjector2_baddress_storage;
assign main_nist_clock_nist_clock_inti_p2_wrdata_en = (main_nist_clock_nist_clock_phaseinjector2_command_issue_re & main_nist_clock_nist_clock_phaseinjector2_command_storage[4]);
assign main_nist_clock_nist_clock_inti_p2_rddata_en = (main_nist_clock_nist_clock_phaseinjector2_command_issue_re & main_nist_clock_nist_clock_phaseinjector2_command_storage[5]);
assign main_nist_clock_nist_clock_inti_p2_wrdata = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage;
assign main_nist_clock_nist_clock_inti_p2_wrdata_mask = 1'd0;

// synthesis translate_off
reg dummy_d_15;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_inti_p3_cas_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p3_cs_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p3_ras_n <= 1'd1;
	main_nist_clock_nist_clock_inti_p3_we_n <= 1'd1;
	if (main_nist_clock_nist_clock_phaseinjector3_command_issue_re) begin
		main_nist_clock_nist_clock_inti_p3_cs_n <= (~main_nist_clock_nist_clock_phaseinjector3_command_storage[0]);
		main_nist_clock_nist_clock_inti_p3_we_n <= (~main_nist_clock_nist_clock_phaseinjector3_command_storage[1]);
		main_nist_clock_nist_clock_inti_p3_cas_n <= (~main_nist_clock_nist_clock_phaseinjector3_command_storage[2]);
		main_nist_clock_nist_clock_inti_p3_ras_n <= (~main_nist_clock_nist_clock_phaseinjector3_command_storage[3]);
	end else begin
		main_nist_clock_nist_clock_inti_p3_cs_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p3_we_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p3_cas_n <= 1'd1;
		main_nist_clock_nist_clock_inti_p3_ras_n <= 1'd1;
	end
// synthesis translate_off
	dummy_d_15 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_inti_p3_address = main_nist_clock_nist_clock_phaseinjector3_address_storage;
assign main_nist_clock_nist_clock_inti_p3_bank = main_nist_clock_nist_clock_phaseinjector3_baddress_storage;
assign main_nist_clock_nist_clock_inti_p3_wrdata_en = (main_nist_clock_nist_clock_phaseinjector3_command_issue_re & main_nist_clock_nist_clock_phaseinjector3_command_storage[4]);
assign main_nist_clock_nist_clock_inti_p3_rddata_en = (main_nist_clock_nist_clock_phaseinjector3_command_issue_re & main_nist_clock_nist_clock_phaseinjector3_command_storage[5]);
assign main_nist_clock_nist_clock_inti_p3_wrdata = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage;
assign main_nist_clock_nist_clock_inti_p3_wrdata_mask = 1'd0;
assign main_nist_clock_nist_clock_sdram_controller_bank0_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset0 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank0_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank1_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset1 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank1_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank2_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset2 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank2_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank3_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset3 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank3_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank4_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset4 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank4_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank5_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset5 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank5_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank6_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset6 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank6_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
assign main_nist_clock_nist_clock_sdram_controller_bank7_open = main_nist_clock_nist_clock_sdram_controller_activate;
assign main_nist_clock_nist_clock_sdram_controller_reset7 = main_nist_clock_nist_clock_sdram_controller_precharge_all;
assign main_nist_clock_nist_clock_sdram_controller_bank7_row0 = main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];

// synthesis translate_off
reg dummy_d_16;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_ce0 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce1 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce2 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce3 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce4 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce5 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce6 <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_ce7 <= 1'd0;
	case (main_nist_clock_nist_clock_sdram_controller_bus_adr[9:7])
		1'd0: begin
			main_nist_clock_nist_clock_sdram_controller_ce0 <= 1'd1;
		end
		1'd1: begin
			main_nist_clock_nist_clock_sdram_controller_ce1 <= 1'd1;
		end
		2'd2: begin
			main_nist_clock_nist_clock_sdram_controller_ce2 <= 1'd1;
		end
		2'd3: begin
			main_nist_clock_nist_clock_sdram_controller_ce3 <= 1'd1;
		end
		3'd4: begin
			main_nist_clock_nist_clock_sdram_controller_ce4 <= 1'd1;
		end
		3'd5: begin
			main_nist_clock_nist_clock_sdram_controller_ce5 <= 1'd1;
		end
		3'd6: begin
			main_nist_clock_nist_clock_sdram_controller_ce6 <= 1'd1;
		end
		3'd7: begin
			main_nist_clock_nist_clock_sdram_controller_ce7 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_16 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sdram_controller_bank_hit = ((((((((main_nist_clock_nist_clock_sdram_controller_bank0_hit & main_nist_clock_nist_clock_sdram_controller_ce0) | (main_nist_clock_nist_clock_sdram_controller_bank1_hit & main_nist_clock_nist_clock_sdram_controller_ce1)) | (main_nist_clock_nist_clock_sdram_controller_bank2_hit & main_nist_clock_nist_clock_sdram_controller_ce2)) | (main_nist_clock_nist_clock_sdram_controller_bank3_hit & main_nist_clock_nist_clock_sdram_controller_ce3)) | (main_nist_clock_nist_clock_sdram_controller_bank4_hit & main_nist_clock_nist_clock_sdram_controller_ce4)) | (main_nist_clock_nist_clock_sdram_controller_bank5_hit & main_nist_clock_nist_clock_sdram_controller_ce5)) | (main_nist_clock_nist_clock_sdram_controller_bank6_hit & main_nist_clock_nist_clock_sdram_controller_ce6)) | (main_nist_clock_nist_clock_sdram_controller_bank7_hit & main_nist_clock_nist_clock_sdram_controller_ce7));
assign main_nist_clock_nist_clock_sdram_controller_bank_idle = ((((((((main_nist_clock_nist_clock_sdram_controller_bank0_idle & main_nist_clock_nist_clock_sdram_controller_ce0) | (main_nist_clock_nist_clock_sdram_controller_bank1_idle & main_nist_clock_nist_clock_sdram_controller_ce1)) | (main_nist_clock_nist_clock_sdram_controller_bank2_idle & main_nist_clock_nist_clock_sdram_controller_ce2)) | (main_nist_clock_nist_clock_sdram_controller_bank3_idle & main_nist_clock_nist_clock_sdram_controller_ce3)) | (main_nist_clock_nist_clock_sdram_controller_bank4_idle & main_nist_clock_nist_clock_sdram_controller_ce4)) | (main_nist_clock_nist_clock_sdram_controller_bank5_idle & main_nist_clock_nist_clock_sdram_controller_ce5)) | (main_nist_clock_nist_clock_sdram_controller_bank6_idle & main_nist_clock_nist_clock_sdram_controller_ce6)) | (main_nist_clock_nist_clock_sdram_controller_bank7_idle & main_nist_clock_nist_clock_sdram_controller_ce7));
assign main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_wait = (~main_nist_clock_nist_clock_sdram_controller_write);
assign main_nist_clock_nist_clock_sdram_controller_refresh_timer_wait = (~main_nist_clock_nist_clock_sdram_controller_refresh);
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_reset_n = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_odt = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_cke = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_cs_n = 1'd0;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p0_bank = main_nist_clock_nist_clock_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_17;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_dfi_p0_address <= 14'd0;
	if (main_nist_clock_nist_clock_sdram_controller_precharge_all) begin
		main_nist_clock_nist_clock_sdram_controller_dfi_p0_address <= 11'd1024;
	end else begin
		if (main_nist_clock_nist_clock_sdram_controller_activate) begin
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_address <= main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
		end else begin
			if ((main_nist_clock_nist_clock_sdram_controller_write | main_nist_clock_nist_clock_sdram_controller_read)) begin
				main_nist_clock_nist_clock_sdram_controller_dfi_p0_address <= {main_nist_clock_nist_clock_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_17 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_reset_n = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_odt = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_cke = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_cs_n = 1'd0;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p1_bank = main_nist_clock_nist_clock_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_18;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_dfi_p1_address <= 14'd0;
	if (main_nist_clock_nist_clock_sdram_controller_precharge_all) begin
		main_nist_clock_nist_clock_sdram_controller_dfi_p1_address <= 11'd1024;
	end else begin
		if (main_nist_clock_nist_clock_sdram_controller_activate) begin
			main_nist_clock_nist_clock_sdram_controller_dfi_p1_address <= main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
		end else begin
			if ((main_nist_clock_nist_clock_sdram_controller_write | main_nist_clock_nist_clock_sdram_controller_read)) begin
				main_nist_clock_nist_clock_sdram_controller_dfi_p1_address <= {main_nist_clock_nist_clock_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_18 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_reset_n = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_odt = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_cke = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_cs_n = 1'd0;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p2_bank = main_nist_clock_nist_clock_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_19;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_dfi_p2_address <= 14'd0;
	if (main_nist_clock_nist_clock_sdram_controller_precharge_all) begin
		main_nist_clock_nist_clock_sdram_controller_dfi_p2_address <= 11'd1024;
	end else begin
		if (main_nist_clock_nist_clock_sdram_controller_activate) begin
			main_nist_clock_nist_clock_sdram_controller_dfi_p2_address <= main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
		end else begin
			if ((main_nist_clock_nist_clock_sdram_controller_write | main_nist_clock_nist_clock_sdram_controller_read)) begin
				main_nist_clock_nist_clock_sdram_controller_dfi_p2_address <= {main_nist_clock_nist_clock_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_19 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_reset_n = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_odt = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_cke = 1'd1;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_cs_n = 1'd0;
assign main_nist_clock_nist_clock_sdram_controller_dfi_p3_bank = main_nist_clock_nist_clock_sdram_controller_bus_adr[9:7];

// synthesis translate_off
reg dummy_d_20;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_dfi_p3_address <= 14'd0;
	if (main_nist_clock_nist_clock_sdram_controller_precharge_all) begin
		main_nist_clock_nist_clock_sdram_controller_dfi_p3_address <= 11'd1024;
	end else begin
		if (main_nist_clock_nist_clock_sdram_controller_activate) begin
			main_nist_clock_nist_clock_sdram_controller_dfi_p3_address <= main_nist_clock_nist_clock_sdram_controller_bus_adr[23:10];
		end else begin
			if ((main_nist_clock_nist_clock_sdram_controller_write | main_nist_clock_nist_clock_sdram_controller_read)) begin
				main_nist_clock_nist_clock_sdram_controller_dfi_p3_address <= {main_nist_clock_nist_clock_sdram_controller_bus_adr[6:0], {3{1'd0}}};
			end
		end
	end
// synthesis translate_off
	dummy_d_20 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sdram_controller_bus_dat_r = {main_nist_clock_nist_clock_sdram_controller_dfi_p3_rddata, main_nist_clock_nist_clock_sdram_controller_dfi_p2_rddata, main_nist_clock_nist_clock_sdram_controller_dfi_p1_rddata, main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata};
assign {main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata, main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata, main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata, main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata} = main_nist_clock_nist_clock_sdram_controller_bus_dat_w;
assign {main_nist_clock_nist_clock_sdram_controller_dfi_p3_wrdata_mask, main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_mask, main_nist_clock_nist_clock_sdram_controller_dfi_p1_wrdata_mask, main_nist_clock_nist_clock_sdram_controller_dfi_p0_wrdata_mask} = (~main_nist_clock_nist_clock_sdram_controller_bus_sel);
assign main_nist_clock_nist_clock_sdram_controller_bank0_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank0_idle) & (main_nist_clock_nist_clock_sdram_controller_bank0_row0 == main_nist_clock_nist_clock_sdram_controller_bank0_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank1_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank1_idle) & (main_nist_clock_nist_clock_sdram_controller_bank1_row0 == main_nist_clock_nist_clock_sdram_controller_bank1_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank2_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank2_idle) & (main_nist_clock_nist_clock_sdram_controller_bank2_row0 == main_nist_clock_nist_clock_sdram_controller_bank2_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank3_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank3_idle) & (main_nist_clock_nist_clock_sdram_controller_bank3_row0 == main_nist_clock_nist_clock_sdram_controller_bank3_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank4_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank4_idle) & (main_nist_clock_nist_clock_sdram_controller_bank4_row0 == main_nist_clock_nist_clock_sdram_controller_bank4_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank5_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank5_idle) & (main_nist_clock_nist_clock_sdram_controller_bank5_row0 == main_nist_clock_nist_clock_sdram_controller_bank5_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank6_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank6_idle) & (main_nist_clock_nist_clock_sdram_controller_bank6_row0 == main_nist_clock_nist_clock_sdram_controller_bank6_row1));
assign main_nist_clock_nist_clock_sdram_controller_bank7_hit = ((~main_nist_clock_nist_clock_sdram_controller_bank7_idle) & (main_nist_clock_nist_clock_sdram_controller_bank7_row0 == main_nist_clock_nist_clock_sdram_controller_bank7_row1));
assign main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_done = (main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count == 1'd0);
assign main_nist_clock_nist_clock_sdram_controller_refresh_timer_done = (main_nist_clock_nist_clock_sdram_controller_refresh_timer_count == 1'd0);

// synthesis translate_off
reg dummy_d_21;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_en <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_dfi_p2_cas_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p2_ras_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p2_we_n <= 1'd1;
	main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_en <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_bus_ack <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_precharge_all <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_activate <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_refresh <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_write <= 1'd0;
	main_nist_clock_nist_clock_sdram_controller_read <= 1'd0;
	builder_minicon_next_state <= 5'd0;
	builder_minicon_next_state <= builder_minicon_state;
	case (builder_minicon_state)
		1'd1: begin
			main_nist_clock_nist_clock_sdram_controller_read <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_en <= 1'd1;
			builder_minicon_next_state <= 2'd2;
		end
		2'd2: begin
			if (main_nist_clock_nist_clock_sdram_controller_dfi_p0_rddata_valid) begin
				main_nist_clock_nist_clock_sdram_controller_bus_ack <= 1'd1;
				builder_minicon_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_nist_clock_nist_clock_sdram_controller_write <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p2_ras_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p2_cas_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p2_we_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p2_wrdata_en <= 1'd1;
			builder_minicon_next_state <= 4'd9;
		end
		3'd4: begin
			main_nist_clock_nist_clock_sdram_controller_bus_ack <= 1'd1;
			builder_minicon_next_state <= 1'd0;
		end
		3'd5: begin
			main_nist_clock_nist_clock_sdram_controller_precharge_all <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd0;
			builder_minicon_next_state <= 4'd14;
		end
		3'd6: begin
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd0;
			builder_minicon_next_state <= 4'd10;
		end
		3'd7: begin
			main_nist_clock_nist_clock_sdram_controller_activate <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd1;
			builder_minicon_next_state <= 4'd12;
		end
		4'd8: begin
			main_nist_clock_nist_clock_sdram_controller_refresh <= 1'd1;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_ras_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_cas_n <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_dfi_p0_we_n <= 1'd1;
			builder_minicon_next_state <= 5'd16;
		end
		4'd9: begin
			builder_minicon_next_state <= 3'd4;
		end
		4'd10: begin
			builder_minicon_next_state <= 4'd11;
		end
		4'd11: begin
			builder_minicon_next_state <= 3'd7;
		end
		4'd12: begin
			builder_minicon_next_state <= 4'd13;
		end
		4'd13: begin
			builder_minicon_next_state <= 1'd0;
		end
		4'd14: begin
			builder_minicon_next_state <= 4'd15;
		end
		4'd15: begin
			builder_minicon_next_state <= 4'd8;
		end
		5'd16: begin
			builder_minicon_next_state <= 5'd17;
		end
		5'd17: begin
			builder_minicon_next_state <= 5'd18;
		end
		5'd18: begin
			builder_minicon_next_state <= 5'd19;
		end
		5'd19: begin
			builder_minicon_next_state <= 5'd20;
		end
		5'd20: begin
			builder_minicon_next_state <= 5'd21;
		end
		5'd21: begin
			builder_minicon_next_state <= 5'd22;
		end
		5'd22: begin
			builder_minicon_next_state <= 5'd23;
		end
		5'd23: begin
			builder_minicon_next_state <= 5'd24;
		end
		5'd24: begin
			builder_minicon_next_state <= 1'd0;
		end
		default: begin
			if (main_nist_clock_nist_clock_sdram_controller_refresh_timer_done) begin
				builder_minicon_next_state <= 3'd5;
			end else begin
				if ((main_nist_clock_nist_clock_sdram_controller_bus_stb & main_nist_clock_nist_clock_sdram_controller_bus_cyc)) begin
					if (main_nist_clock_nist_clock_sdram_controller_bank_hit) begin
						if (main_nist_clock_nist_clock_sdram_controller_bus_we) begin
							builder_minicon_next_state <= 2'd3;
						end else begin
							builder_minicon_next_state <= 1'd1;
						end
					end else begin
						if ((~main_nist_clock_nist_clock_sdram_controller_bank_idle)) begin
							if (main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_done) begin
								builder_minicon_next_state <= 3'd6;
							end
						end else begin
							builder_minicon_next_state <= 3'd7;
						end
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_21 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_data_port_adr = main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[14:4];

// synthesis translate_off
reg dummy_d_22;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_data_port_we <= 64'd0;
	main_nist_clock_nist_clock_data_port_dat_w <= 512'd0;
	if (main_nist_clock_nist_clock_write_from_slave) begin
		main_nist_clock_nist_clock_data_port_dat_w <= main_nist_clock_nist_clock_bridge_if_bus_dat_r;
		main_nist_clock_nist_clock_data_port_we <= {64{1'd1}};
	end else begin
		main_nist_clock_nist_clock_data_port_dat_w <= {16{main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_w}};
		if ((((main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cyc & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_stb) & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_we) & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack)) begin
			main_nist_clock_nist_clock_data_port_we <= {({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 1'd0)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 1'd1)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 2'd2)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 2'd3)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 3'd4)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 3'd5)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 3'd6)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 3'd7)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd8)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd9)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd10)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd11)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd12)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd13)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd14)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel), ({4{(main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0] == 4'd15)}} & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel)};
		end
	end
// synthesis translate_off
	dummy_d_22 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_bridge_if_bus_dat_w = main_nist_clock_nist_clock_data_port_dat_r;
assign main_nist_clock_nist_clock_bridge_if_bus_sel = 64'd18446744073709551615;

// synthesis translate_off
reg dummy_d_23;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= 32'd0;
	case (main_nist_clock_nist_clock_adr_offset_r)
		1'd0: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[511:480];
		end
		1'd1: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[479:448];
		end
		2'd2: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[447:416];
		end
		2'd3: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[415:384];
		end
		3'd4: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[383:352];
		end
		3'd5: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[351:320];
		end
		3'd6: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[319:288];
		end
		3'd7: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[287:256];
		end
		4'd8: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[255:224];
		end
		4'd9: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[223:192];
		end
		4'd10: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[191:160];
		end
		4'd11: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[159:128];
		end
		4'd12: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[127:96];
		end
		4'd13: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[95:64];
		end
		4'd14: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[63:32];
		end
		default: begin
			main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r <= main_nist_clock_nist_clock_data_port_dat_r[31:0];
		end
	endcase
// synthesis translate_off
	dummy_d_23 <= dummy_s;
// synthesis translate_on
end
assign {main_nist_clock_nist_clock_tag_do_dirty, main_nist_clock_nist_clock_tag_do_tag} = main_nist_clock_nist_clock_tag_port_dat_r;
assign main_nist_clock_nist_clock_tag_port_dat_w = {main_nist_clock_nist_clock_tag_di_dirty, main_nist_clock_nist_clock_tag_di_tag};
assign main_nist_clock_nist_clock_tag_port_adr = main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[14:4];
assign main_nist_clock_nist_clock_tag_di_tag = main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[29:15];
assign main_nist_clock_nist_clock_bridge_if_bus_adr = {main_nist_clock_nist_clock_tag_do_tag, main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[14:4]};

// synthesis translate_off
reg dummy_d_24;
// synthesis translate_on
always @(*) begin
	main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack <= 1'd0;
	main_nist_clock_nist_clock_bridge_if_bus_cyc <= 1'd0;
	main_nist_clock_nist_clock_bridge_if_bus_stb <= 1'd0;
	main_nist_clock_nist_clock_bridge_if_bus_we <= 1'd0;
	main_nist_clock_nist_clock_write_from_slave <= 1'd0;
	main_nist_clock_nist_clock_tag_port_we <= 1'd0;
	main_nist_clock_nist_clock_tag_di_dirty <= 1'd0;
	main_nist_clock_nist_clock_word_clr <= 1'd0;
	main_nist_clock_nist_clock_word_inc <= 1'd0;
	builder_fullmemorywe_next_state <= 3'd0;
	builder_fullmemorywe_next_state <= builder_fullmemorywe_state;
	case (builder_fullmemorywe_state)
		1'd1: begin
			main_nist_clock_nist_clock_word_clr <= 1'd1;
			if ((main_nist_clock_nist_clock_tag_do_tag == main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[29:15])) begin
				main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack <= 1'd1;
				if (main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_we) begin
					main_nist_clock_nist_clock_tag_di_dirty <= 1'd1;
					main_nist_clock_nist_clock_tag_port_we <= 1'd1;
				end
				builder_fullmemorywe_next_state <= 1'd0;
			end else begin
				if (main_nist_clock_nist_clock_tag_do_dirty) begin
					builder_fullmemorywe_next_state <= 2'd2;
				end else begin
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			main_nist_clock_nist_clock_bridge_if_bus_stb <= 1'd1;
			main_nist_clock_nist_clock_bridge_if_bus_cyc <= 1'd1;
			main_nist_clock_nist_clock_bridge_if_bus_we <= 1'd1;
			if (main_nist_clock_nist_clock_bridge_if_bus_ack) begin
				main_nist_clock_nist_clock_word_inc <= 1'd1;
				if (1'd1) begin
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			main_nist_clock_nist_clock_tag_port_we <= 1'd1;
			main_nist_clock_nist_clock_word_clr <= 1'd1;
			builder_fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			main_nist_clock_nist_clock_bridge_if_bus_stb <= 1'd1;
			main_nist_clock_nist_clock_bridge_if_bus_cyc <= 1'd1;
			main_nist_clock_nist_clock_bridge_if_bus_we <= 1'd0;
			if (main_nist_clock_nist_clock_bridge_if_bus_ack) begin
				main_nist_clock_nist_clock_write_from_slave <= 1'd1;
				main_nist_clock_nist_clock_word_inc <= 1'd1;
				if (1'd1) begin
					builder_fullmemorywe_next_state <= 1'd1;
				end else begin
					builder_fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cyc & main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_stb)) begin
				builder_fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_24 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_spiflash_bus_dat_r = main_nist_clock_spiflash_sr;

// synthesis translate_off
reg dummy_d_25;
// synthesis translate_on
always @(*) begin
	spiflash_cs_n <= 1'd1;
	main_nist_clock_clk <= 1'd0;
	main_nist_clock_spiflash_status <= 1'd0;
	main_nist_clock_spiflash_o <= 4'd0;
	main_nist_clock_spiflash_oe <= 1'd0;
	if (main_nist_clock_spiflash_bitbang_en_storage) begin
		main_nist_clock_clk <= main_nist_clock_spiflash_bitbang_storage[1];
		spiflash_cs_n <= main_nist_clock_spiflash_bitbang_storage[2];
		if (main_nist_clock_spiflash_bitbang_storage[3]) begin
			main_nist_clock_spiflash_oe <= 1'd0;
		end else begin
			main_nist_clock_spiflash_oe <= 1'd1;
		end
		if (main_nist_clock_spiflash_bitbang_storage[1]) begin
			main_nist_clock_spiflash_status <= main_nist_clock_spiflash_i0[1];
		end
		main_nist_clock_spiflash_o <= {{3{1'd1}}, main_nist_clock_spiflash_bitbang_storage[0]};
	end else begin
		main_nist_clock_clk <= main_nist_clock_spiflash_clk;
		spiflash_cs_n <= main_nist_clock_spiflash_cs_n1;
		main_nist_clock_spiflash_o <= main_nist_clock_spiflash_sr[31:28];
		main_nist_clock_spiflash_oe <= main_nist_clock_spiflash_dq_oe;
	end
// synthesis translate_off
	dummy_d_25 <= dummy_s;
// synthesis translate_on
end
assign main_ethphy_mode_status = main_ethphy_mode0;
assign main_ethphy_eth_tick = (main_ethphy_eth_counter == 1'd0);
assign main_ethphy_i = main_ethphy_eth_tick;
assign main_ethphy_sys_tick = main_ethphy_o;
assign main_ethphy_o = (main_ethphy_toggle_o ^ main_ethphy_toggle_o_r);

// synthesis translate_off
reg dummy_d_26;
// synthesis translate_on
always @(*) begin
	main_ethphy_mode1 <= 1'd0;
	main_ethphy_update_mode <= 1'd0;
	main_ethphy_sys_counter_reset <= 1'd0;
	main_ethphy_sys_counter_ce <= 1'd0;
	builder_liteethphygmiimii_next_state <= 2'd0;
	builder_liteethphygmiimii_next_state <= builder_liteethphygmiimii_state;
	case (builder_liteethphygmiimii_state)
		1'd1: begin
			main_ethphy_sys_counter_ce <= 1'd1;
			if (main_ethphy_sys_tick) begin
				builder_liteethphygmiimii_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_ethphy_update_mode <= 1'd1;
			if ((main_ethphy_sys_counter > 11'd1075)) begin
				main_ethphy_mode1 <= 1'd1;
			end else begin
				main_ethphy_mode1 <= 1'd0;
			end
			builder_liteethphygmiimii_next_state <= 1'd0;
		end
		default: begin
			main_ethphy_sys_counter_reset <= 1'd1;
			if (main_ethphy_sys_tick) begin
				builder_liteethphygmiimii_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_26 <= dummy_s;
// synthesis translate_on
end
assign eth_rx_clk = eth_clocks_rx;
assign eth_rst_n = (~main_ethphy_storage);
assign main_ethphy_liteethphygmiimiitx_demux_sel = (main_ethphy_mode0 == 1'd1);
assign main_ethphy_liteethphygmiimiitx_demux_sink_stb = main_ethphy_liteethphygmiimiitx_sink_sink_stb0;
assign main_ethphy_liteethphygmiimiitx_sink_sink_ack0 = main_ethphy_liteethphygmiimiitx_demux_sink_ack;
assign main_ethphy_liteethphygmiimiitx_demux_sink_eop = main_ethphy_liteethphygmiimiitx_sink_sink_eop0;
assign main_ethphy_liteethphygmiimiitx_demux_sink_payload_data = main_ethphy_liteethphygmiimiitx_sink_sink_payload_data0;
assign main_ethphy_liteethphygmiimiitx_demux_sink_payload_last_be = main_ethphy_liteethphygmiimiitx_sink_sink_payload_last_be0;
assign main_ethphy_liteethphygmiimiitx_demux_sink_payload_error = main_ethphy_liteethphygmiimiitx_sink_sink_payload_error0;
assign main_ethphy_liteethphygmiimiitx_gmii_tx_sink_stb = main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_stb;
assign main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_ack = main_ethphy_liteethphygmiimiitx_gmii_tx_sink_ack;
assign main_ethphy_liteethphygmiimiitx_gmii_tx_sink_eop = main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_eop;
assign main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_data = main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_data;
assign main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_last_be = main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_last_be;
assign main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_error = main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_error;
assign main_ethphy_liteethphygmiimiitx_sink_sink_stb1 = main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_stb;
assign main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_ack = main_ethphy_liteethphygmiimiitx_sink_sink_ack1;
assign main_ethphy_liteethphygmiimiitx_sink_sink_eop1 = main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_eop;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_data1 = main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_data;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_last_be1 = main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_last_be;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_error1 = main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_error;
assign eth_tx_er = 1'd0;
assign main_ethphy_liteethphygmiimiitx_converter_sink_stb = main_ethphy_liteethphygmiimiitx_sink_sink_stb1;
assign main_ethphy_liteethphygmiimiitx_converter_sink_payload_data = main_ethphy_liteethphygmiimiitx_sink_sink_payload_data1;
assign main_ethphy_liteethphygmiimiitx_sink_sink_ack1 = main_ethphy_liteethphygmiimiitx_converter_sink_ack;
assign main_ethphy_liteethphygmiimiitx_converter_source_ack = 1'd1;
assign main_ethphy_liteethphygmiimiitx_converter_last = (main_ethphy_liteethphygmiimiitx_converter_mux == 1'd1);
assign main_ethphy_liteethphygmiimiitx_converter_source_stb = main_ethphy_liteethphygmiimiitx_converter_sink_stb;
assign main_ethphy_liteethphygmiimiitx_converter_source_eop = (main_ethphy_liteethphygmiimiitx_converter_sink_eop & main_ethphy_liteethphygmiimiitx_converter_last);
assign main_ethphy_liteethphygmiimiitx_converter_sink_ack = (main_ethphy_liteethphygmiimiitx_converter_last & main_ethphy_liteethphygmiimiitx_converter_source_ack);

// synthesis translate_off
reg dummy_d_27;
// synthesis translate_on
always @(*) begin
	main_ethphy_liteethphygmiimiitx_converter_source_payload_data <= 4'd0;
	case (main_ethphy_liteethphygmiimiitx_converter_mux)
		1'd0: begin
			main_ethphy_liteethphygmiimiitx_converter_source_payload_data <= main_ethphy_liteethphygmiimiitx_converter_sink_payload_data[3:0];
		end
		default: begin
			main_ethphy_liteethphygmiimiitx_converter_source_payload_data <= main_ethphy_liteethphygmiimiitx_converter_sink_payload_data[7:4];
		end
	endcase
// synthesis translate_off
	dummy_d_27 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_28;
// synthesis translate_on
always @(*) begin
	main_ethphy_liteethphygmiimiitx_demux_sink_ack <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_stb <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_eop <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_data <= 8'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_last_be <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_error <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_stb <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_eop <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_data <= 8'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_last_be <= 1'd0;
	main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_error <= 1'd0;
	case (main_ethphy_liteethphygmiimiitx_demux_sel)
		1'd0: begin
			main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_stb <= main_ethphy_liteethphygmiimiitx_demux_sink_stb;
			main_ethphy_liteethphygmiimiitx_demux_sink_ack <= main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_ack;
			main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_eop <= main_ethphy_liteethphygmiimiitx_demux_sink_eop;
			main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_data <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_data;
			main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_last_be <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_last_be;
			main_ethphy_liteethphygmiimiitx_demux_endpoint0_source_payload_error <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_error;
		end
		1'd1: begin
			main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_stb <= main_ethphy_liteethphygmiimiitx_demux_sink_stb;
			main_ethphy_liteethphygmiimiitx_demux_sink_ack <= main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_ack;
			main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_eop <= main_ethphy_liteethphygmiimiitx_demux_sink_eop;
			main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_data <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_data;
			main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_last_be <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_last_be;
			main_ethphy_liteethphygmiimiitx_demux_endpoint1_source_payload_error <= main_ethphy_liteethphygmiimiitx_demux_sink_payload_error;
		end
	endcase
// synthesis translate_off
	dummy_d_28 <= dummy_s;
// synthesis translate_on
end
assign main_ethphy_liteethphygmiimiirx_mux_sel = (main_ethphy_mode0 == 1'd1);
assign main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_stb = main_ethphy_liteethphygmiimiirx_gmii_rx_source_stb;
assign main_ethphy_liteethphygmiimiirx_gmii_rx_source_ack = main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_ack;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_eop = main_ethphy_liteethphygmiimiirx_gmii_rx_source_eop;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_data = main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_data;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_last_be = main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_last_be;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_error = main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_error;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_stb = main_ethphy_liteethphygmiimiirx_source_source_stb1;
assign main_ethphy_liteethphygmiimiirx_source_source_ack1 = main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_ack;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_eop = main_ethphy_liteethphygmiimiirx_source_source_eop1;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_data = main_ethphy_liteethphygmiimiirx_source_source_payload_data1;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_last_be = main_ethphy_liteethphygmiimiirx_source_source_payload_last_be1;
assign main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_error = main_ethphy_liteethphygmiimiirx_source_source_payload_error1;
assign main_ethphy_liteethphygmiimiirx_source_source_stb0 = main_ethphy_liteethphygmiimiirx_mux_source_stb;
assign main_ethphy_liteethphygmiimiirx_mux_source_ack = main_ethphy_liteethphygmiimiirx_source_source_ack0;
assign main_ethphy_liteethphygmiimiirx_source_source_eop0 = main_ethphy_liteethphygmiimiirx_mux_source_eop;
assign main_ethphy_liteethphygmiimiirx_source_source_payload_data0 = main_ethphy_liteethphygmiimiirx_mux_source_payload_data;
assign main_ethphy_liteethphygmiimiirx_source_source_payload_last_be0 = main_ethphy_liteethphygmiimiirx_mux_source_payload_last_be;
assign main_ethphy_liteethphygmiimiirx_source_source_payload_error0 = main_ethphy_liteethphygmiimiirx_mux_source_payload_error;
assign main_ethphy_liteethphygmiimiirx_gmii_rx_source_eop = ((~main_ethphy_liteethphygmiimiirx_pads_d_rx_dv) & main_ethphy_liteethphygmiimiirx_gmii_rx_rx_dv_d);
assign main_ethphy_liteethphygmiimiirx_converter_sink_eop = (~main_ethphy_liteethphygmiimiirx_pads_d_rx_dv);
assign main_ethphy_liteethphygmiimiirx_source_source_stb1 = main_ethphy_liteethphygmiimiirx_converter_source_stb;
assign main_ethphy_liteethphygmiimiirx_converter_source_ack = main_ethphy_liteethphygmiimiirx_source_source_ack1;
assign main_ethphy_liteethphygmiimiirx_source_source_eop1 = main_ethphy_liteethphygmiimiirx_converter_source_eop;
assign main_ethphy_liteethphygmiimiirx_source_source_payload_data1 = main_ethphy_liteethphygmiimiirx_converter_source_payload_data;
assign main_ethphy_liteethphygmiimiirx_converter_sink_ack = ((~main_ethphy_liteethphygmiimiirx_converter_strobe_all) | main_ethphy_liteethphygmiimiirx_converter_source_ack);
assign main_ethphy_liteethphygmiimiirx_converter_source_stb = main_ethphy_liteethphygmiimiirx_converter_strobe_all;
assign main_ethphy_liteethphygmiimiirx_converter_load_part = (main_ethphy_liteethphygmiimiirx_converter_sink_stb & main_ethphy_liteethphygmiimiirx_converter_sink_ack);

// synthesis translate_off
reg dummy_d_29;
// synthesis translate_on
always @(*) begin
	main_ethphy_liteethphygmiimiirx_mux_source_stb <= 1'd0;
	main_ethphy_liteethphygmiimiirx_mux_source_eop <= 1'd0;
	main_ethphy_liteethphygmiimiirx_mux_source_payload_data <= 8'd0;
	main_ethphy_liteethphygmiimiirx_mux_source_payload_last_be <= 1'd0;
	main_ethphy_liteethphygmiimiirx_mux_source_payload_error <= 1'd0;
	main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_ack <= 1'd0;
	main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_ack <= 1'd0;
	case (main_ethphy_liteethphygmiimiirx_mux_sel)
		1'd0: begin
			main_ethphy_liteethphygmiimiirx_mux_source_stb <= main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_stb;
			main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_ack <= main_ethphy_liteethphygmiimiirx_mux_source_ack;
			main_ethphy_liteethphygmiimiirx_mux_source_eop <= main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_eop;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_data <= main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_data;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_last_be <= main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_last_be;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_error <= main_ethphy_liteethphygmiimiirx_mux_endpoint0_sink_payload_error;
		end
		1'd1: begin
			main_ethphy_liteethphygmiimiirx_mux_source_stb <= main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_stb;
			main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_ack <= main_ethphy_liteethphygmiimiirx_mux_source_ack;
			main_ethphy_liteethphygmiimiirx_mux_source_eop <= main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_eop;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_data <= main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_data;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_last_be <= main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_last_be;
			main_ethphy_liteethphygmiimiirx_mux_source_payload_error <= main_ethphy_liteethphygmiimiirx_mux_endpoint1_sink_payload_error;
		end
	endcase
// synthesis translate_off
	dummy_d_29 <= dummy_s;
// synthesis translate_on
end
assign main_tx_cdc_sink_stb = main_source_stb;
assign main_source_ack = main_tx_cdc_sink_ack;
assign main_tx_cdc_sink_eop = main_source_eop;
assign main_tx_cdc_sink_payload_data = main_source_payload_data;
assign main_tx_cdc_sink_payload_last_be = main_source_payload_last_be;
assign main_tx_cdc_sink_payload_error = main_source_payload_error;
assign main_sink_stb = main_rx_cdc_source_stb;
assign main_rx_cdc_source_ack = main_sink_ack;
assign main_sink_eop = main_rx_cdc_source_eop;
assign main_sink_payload_data = main_rx_cdc_source_payload_data;
assign main_sink_payload_last_be = main_rx_cdc_source_payload_last_be;
assign main_sink_payload_error = main_rx_cdc_source_payload_error;
assign main_ps_preamble_error_i = main_preamble_checker_error;
assign main_ps_crc_error_i = main_crc32_checker_error;
assign main_tx_converter_sink_sink_stb = main_tx_cdc_source_stb;
assign main_tx_cdc_source_ack = main_tx_converter_sink_sink_ack;
assign main_tx_converter_sink_sink_eop = main_tx_cdc_source_eop;
assign main_tx_converter_sink_sink_payload_data = main_tx_cdc_source_payload_data;
assign main_tx_converter_sink_sink_payload_last_be = main_tx_cdc_source_payload_last_be;
assign main_tx_converter_sink_sink_payload_error = main_tx_cdc_source_payload_error;
assign main_tx_last_be_sink_stb = main_tx_converter_source_source_stb;
assign main_tx_converter_source_source_ack = main_tx_last_be_sink_ack;
assign main_tx_last_be_sink_eop = main_tx_converter_source_source_eop;
assign main_tx_last_be_sink_payload_data = main_tx_converter_source_source_payload_data;
assign main_tx_last_be_sink_payload_last_be = main_tx_converter_source_source_payload_last_be;
assign main_tx_last_be_sink_payload_error = main_tx_converter_source_source_payload_error;
assign main_padding_inserter_sink_stb = main_tx_last_be_source_stb;
assign main_tx_last_be_source_ack = main_padding_inserter_sink_ack;
assign main_padding_inserter_sink_eop = main_tx_last_be_source_eop;
assign main_padding_inserter_sink_payload_data = main_tx_last_be_source_payload_data;
assign main_padding_inserter_sink_payload_last_be = main_tx_last_be_source_payload_last_be;
assign main_padding_inserter_sink_payload_error = main_tx_last_be_source_payload_error;
assign main_crc32_inserter_sink_stb = main_padding_inserter_source_stb;
assign main_padding_inserter_source_ack = main_crc32_inserter_sink_ack;
assign main_crc32_inserter_sink_eop = main_padding_inserter_source_eop;
assign main_crc32_inserter_sink_payload_data = main_padding_inserter_source_payload_data;
assign main_crc32_inserter_sink_payload_last_be = main_padding_inserter_source_payload_last_be;
assign main_crc32_inserter_sink_payload_error = main_padding_inserter_source_payload_error;
assign main_preamble_inserter_sink_stb = main_crc32_inserter_source_stb;
assign main_crc32_inserter_source_ack = main_preamble_inserter_sink_ack;
assign main_preamble_inserter_sink_eop = main_crc32_inserter_source_eop;
assign main_preamble_inserter_sink_payload_data = main_crc32_inserter_source_payload_data;
assign main_preamble_inserter_sink_payload_last_be = main_crc32_inserter_source_payload_last_be;
assign main_preamble_inserter_sink_payload_error = main_crc32_inserter_source_payload_error;
assign main_tx_gap_inserter_sink_stb = main_preamble_inserter_source_stb;
assign main_preamble_inserter_source_ack = main_tx_gap_inserter_sink_ack;
assign main_tx_gap_inserter_sink_eop = main_preamble_inserter_source_eop;
assign main_tx_gap_inserter_sink_payload_data = main_preamble_inserter_source_payload_data;
assign main_tx_gap_inserter_sink_payload_last_be = main_preamble_inserter_source_payload_last_be;
assign main_tx_gap_inserter_sink_payload_error = main_preamble_inserter_source_payload_error;
assign main_ethphy_liteethphygmiimiitx_sink_sink_stb0 = main_tx_gap_inserter_source_stb;
assign main_tx_gap_inserter_source_ack = main_ethphy_liteethphygmiimiitx_sink_sink_ack0;
assign main_ethphy_liteethphygmiimiitx_sink_sink_eop0 = main_tx_gap_inserter_source_eop;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_data0 = main_tx_gap_inserter_source_payload_data;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_last_be0 = main_tx_gap_inserter_source_payload_last_be;
assign main_ethphy_liteethphygmiimiitx_sink_sink_payload_error0 = main_tx_gap_inserter_source_payload_error;
assign main_preamble_checker_sink_stb = main_ethphy_liteethphygmiimiirx_source_source_stb0;
assign main_ethphy_liteethphygmiimiirx_source_source_ack0 = main_preamble_checker_sink_ack;
assign main_preamble_checker_sink_eop = main_ethphy_liteethphygmiimiirx_source_source_eop0;
assign main_preamble_checker_sink_payload_data = main_ethphy_liteethphygmiimiirx_source_source_payload_data0;
assign main_preamble_checker_sink_payload_last_be = main_ethphy_liteethphygmiimiirx_source_source_payload_last_be0;
assign main_preamble_checker_sink_payload_error = main_ethphy_liteethphygmiimiirx_source_source_payload_error0;
assign main_crc32_checker_sink_sink_stb = main_preamble_checker_source_stb;
assign main_preamble_checker_source_ack = main_crc32_checker_sink_sink_ack;
assign main_crc32_checker_sink_sink_eop = main_preamble_checker_source_eop;
assign main_crc32_checker_sink_sink_payload_data = main_preamble_checker_source_payload_data;
assign main_crc32_checker_sink_sink_payload_last_be = main_preamble_checker_source_payload_last_be;
assign main_crc32_checker_sink_sink_payload_error = main_preamble_checker_source_payload_error;
assign main_padding_checker_sink_stb = main_crc32_checker_source_source_stb;
assign main_crc32_checker_source_source_ack = main_padding_checker_sink_ack;
assign main_padding_checker_sink_eop = main_crc32_checker_source_source_eop;
assign main_padding_checker_sink_payload_data = main_crc32_checker_source_source_payload_data;
assign main_padding_checker_sink_payload_last_be = main_crc32_checker_source_source_payload_last_be;
assign main_padding_checker_sink_payload_error = main_crc32_checker_source_source_payload_error;
assign main_rx_last_be_sink_stb = main_padding_checker_source_stb;
assign main_padding_checker_source_ack = main_rx_last_be_sink_ack;
assign main_rx_last_be_sink_eop = main_padding_checker_source_eop;
assign main_rx_last_be_sink_payload_data = main_padding_checker_source_payload_data;
assign main_rx_last_be_sink_payload_last_be = main_padding_checker_source_payload_last_be;
assign main_rx_last_be_sink_payload_error = main_padding_checker_source_payload_error;
assign main_rx_converter_sink_sink_stb = main_rx_last_be_source_stb;
assign main_rx_last_be_source_ack = main_rx_converter_sink_sink_ack;
assign main_rx_converter_sink_sink_eop = main_rx_last_be_source_eop;
assign main_rx_converter_sink_sink_payload_data = main_rx_last_be_source_payload_data;
assign main_rx_converter_sink_sink_payload_last_be = main_rx_last_be_source_payload_last_be;
assign main_rx_converter_sink_sink_payload_error = main_rx_last_be_source_payload_error;
assign main_rx_cdc_sink_stb = main_rx_converter_source_source_stb;
assign main_rx_converter_source_source_ack = main_rx_cdc_sink_ack;
assign main_rx_cdc_sink_eop = main_rx_converter_source_source_eop;
assign main_rx_cdc_sink_payload_data = main_rx_converter_source_source_payload_data;
assign main_rx_cdc_sink_payload_last_be = main_rx_converter_source_source_payload_last_be;
assign main_rx_cdc_sink_payload_error = main_rx_converter_source_source_payload_error;

// synthesis translate_off
reg dummy_d_30;
// synthesis translate_on
always @(*) begin
	main_tx_gap_inserter_sink_ack <= 1'd0;
	main_tx_gap_inserter_source_stb <= 1'd0;
	main_tx_gap_inserter_source_eop <= 1'd0;
	main_tx_gap_inserter_source_payload_data <= 8'd0;
	main_tx_gap_inserter_source_payload_last_be <= 1'd0;
	main_tx_gap_inserter_source_payload_error <= 1'd0;
	main_tx_gap_inserter_counter_reset <= 1'd0;
	main_tx_gap_inserter_counter_ce <= 1'd0;
	builder_liteethmacgap_next_state <= 1'd0;
	builder_liteethmacgap_next_state <= builder_liteethmacgap_state;
	case (builder_liteethmacgap_state)
		1'd1: begin
			main_tx_gap_inserter_counter_ce <= 1'd1;
			if ((main_tx_gap_inserter_counter == 4'd11)) begin
				builder_liteethmacgap_next_state <= 1'd0;
			end
		end
		default: begin
			main_tx_gap_inserter_counter_reset <= 1'd1;
			main_tx_gap_inserter_source_stb <= main_tx_gap_inserter_sink_stb;
			main_tx_gap_inserter_sink_ack <= main_tx_gap_inserter_source_ack;
			main_tx_gap_inserter_source_eop <= main_tx_gap_inserter_sink_eop;
			main_tx_gap_inserter_source_payload_data <= main_tx_gap_inserter_sink_payload_data;
			main_tx_gap_inserter_source_payload_last_be <= main_tx_gap_inserter_sink_payload_last_be;
			main_tx_gap_inserter_source_payload_error <= main_tx_gap_inserter_sink_payload_error;
			if (((main_tx_gap_inserter_sink_stb & main_tx_gap_inserter_sink_eop) & main_tx_gap_inserter_sink_ack)) begin
				builder_liteethmacgap_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_30 <= dummy_s;
// synthesis translate_on
end
assign main_preamble_inserter_source_payload_last_be = main_preamble_inserter_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_31;
// synthesis translate_on
always @(*) begin
	main_preamble_inserter_sink_ack <= 1'd0;
	main_preamble_inserter_source_stb <= 1'd0;
	main_preamble_inserter_source_eop <= 1'd0;
	main_preamble_inserter_source_payload_data <= 8'd0;
	main_preamble_inserter_source_payload_error <= 1'd0;
	main_preamble_inserter_clr_cnt <= 1'd0;
	main_preamble_inserter_inc_cnt <= 1'd0;
	builder_liteethmacpreambleinserter_next_state <= 2'd0;
	main_preamble_inserter_source_payload_data <= main_preamble_inserter_sink_payload_data;
	builder_liteethmacpreambleinserter_next_state <= builder_liteethmacpreambleinserter_state;
	case (builder_liteethmacpreambleinserter_state)
		1'd1: begin
			main_preamble_inserter_source_stb <= 1'd1;
			case (main_preamble_inserter_cnt)
				1'd0: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[55:48];
				end
				default: begin
					main_preamble_inserter_source_payload_data <= main_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((main_preamble_inserter_cnt == 3'd7)) begin
				if (main_preamble_inserter_source_ack) begin
					builder_liteethmacpreambleinserter_next_state <= 2'd2;
				end
			end else begin
				main_preamble_inserter_inc_cnt <= main_preamble_inserter_source_ack;
			end
		end
		2'd2: begin
			main_preamble_inserter_source_stb <= main_preamble_inserter_sink_stb;
			main_preamble_inserter_sink_ack <= main_preamble_inserter_source_ack;
			main_preamble_inserter_source_eop <= main_preamble_inserter_sink_eop;
			main_preamble_inserter_source_payload_error <= main_preamble_inserter_sink_payload_error;
			if (((main_preamble_inserter_sink_stb & main_preamble_inserter_sink_eop) & main_preamble_inserter_source_ack)) begin
				builder_liteethmacpreambleinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_preamble_inserter_sink_ack <= 1'd1;
			main_preamble_inserter_clr_cnt <= 1'd1;
			if (main_preamble_inserter_sink_stb) begin
				main_preamble_inserter_sink_ack <= 1'd0;
				builder_liteethmacpreambleinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_31 <= dummy_s;
// synthesis translate_on
end
assign main_preamble_checker_source_payload_data = main_preamble_checker_sink_payload_data;
assign main_preamble_checker_source_payload_last_be = main_preamble_checker_sink_payload_last_be;

// synthesis translate_off
reg dummy_d_32;
// synthesis translate_on
always @(*) begin
	main_preamble_checker_sink_ack <= 1'd0;
	main_preamble_checker_source_stb <= 1'd0;
	main_preamble_checker_source_eop <= 1'd0;
	main_preamble_checker_source_payload_error <= 1'd0;
	main_preamble_checker_error <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= 1'd0;
	builder_liteethmacpreamblechecker_next_state <= builder_liteethmacpreamblechecker_state;
	case (builder_liteethmacpreamblechecker_state)
		1'd1: begin
			main_preamble_checker_source_stb <= main_preamble_checker_sink_stb;
			main_preamble_checker_sink_ack <= main_preamble_checker_source_ack;
			main_preamble_checker_source_eop <= main_preamble_checker_sink_eop;
			main_preamble_checker_source_payload_error <= main_preamble_checker_sink_payload_error;
			if (((main_preamble_checker_source_stb & main_preamble_checker_source_eop) & main_preamble_checker_source_ack)) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd0;
			end
		end
		default: begin
			main_preamble_checker_sink_ack <= 1'd1;
			if (((main_preamble_checker_sink_stb & (~main_preamble_checker_sink_eop)) & (main_preamble_checker_sink_payload_data == 8'd213))) begin
				builder_liteethmacpreamblechecker_next_state <= 1'd1;
			end
			if ((main_preamble_checker_sink_stb & main_preamble_checker_sink_eop)) begin
				main_preamble_checker_error <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_32 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_inserter_cnt_done = (main_crc32_inserter_cnt == 1'd0);
assign main_crc32_inserter_data1 = main_crc32_inserter_data0;
assign main_crc32_inserter_last = main_crc32_inserter_reg;
assign main_crc32_inserter_value = (~{main_crc32_inserter_reg[0], main_crc32_inserter_reg[1], main_crc32_inserter_reg[2], main_crc32_inserter_reg[3], main_crc32_inserter_reg[4], main_crc32_inserter_reg[5], main_crc32_inserter_reg[6], main_crc32_inserter_reg[7], main_crc32_inserter_reg[8], main_crc32_inserter_reg[9], main_crc32_inserter_reg[10], main_crc32_inserter_reg[11], main_crc32_inserter_reg[12], main_crc32_inserter_reg[13], main_crc32_inserter_reg[14], main_crc32_inserter_reg[15], main_crc32_inserter_reg[16], main_crc32_inserter_reg[17], main_crc32_inserter_reg[18], main_crc32_inserter_reg[19], main_crc32_inserter_reg[20], main_crc32_inserter_reg[21], main_crc32_inserter_reg[22], main_crc32_inserter_reg[23], main_crc32_inserter_reg[24], main_crc32_inserter_reg[25], main_crc32_inserter_reg[26], main_crc32_inserter_reg[27], main_crc32_inserter_reg[28], main_crc32_inserter_reg[29], main_crc32_inserter_reg[30], main_crc32_inserter_reg[31]});
assign main_crc32_inserter_error = (main_crc32_inserter_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_33;
// synthesis translate_on
always @(*) begin
	main_crc32_inserter_next <= 32'd0;
	main_crc32_inserter_next[0] <= (((main_crc32_inserter_last[24] ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[1] <= (((((((main_crc32_inserter_last[25] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[2] <= (((((((((main_crc32_inserter_last[26] ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[3] <= (((((((main_crc32_inserter_last[27] ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[4] <= (((((((((main_crc32_inserter_last[28] ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[5] <= (((((((((((((main_crc32_inserter_last[29] ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[6] <= (((((((((((main_crc32_inserter_last[30] ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[7] <= (((((((((main_crc32_inserter_last[31] ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[8] <= ((((((((main_crc32_inserter_last[0] ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[9] <= ((((((((main_crc32_inserter_last[1] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[10] <= ((((((((main_crc32_inserter_last[2] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[11] <= ((((((((main_crc32_inserter_last[3] ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[12] <= ((((((((((((main_crc32_inserter_last[4] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[13] <= ((((((((((((main_crc32_inserter_last[5] ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[14] <= ((((((((((main_crc32_inserter_last[6] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]);
	main_crc32_inserter_next[15] <= ((((((((main_crc32_inserter_last[7] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]);
	main_crc32_inserter_next[16] <= ((((((main_crc32_inserter_last[8] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[17] <= ((((((main_crc32_inserter_last[9] ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[18] <= ((((((main_crc32_inserter_last[10] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]);
	main_crc32_inserter_next[19] <= ((((main_crc32_inserter_last[11] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]);
	main_crc32_inserter_next[20] <= ((main_crc32_inserter_last[12] ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]);
	main_crc32_inserter_next[21] <= ((main_crc32_inserter_last[13] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]);
	main_crc32_inserter_next[22] <= ((main_crc32_inserter_last[14] ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[23] <= ((((((main_crc32_inserter_last[15] ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_data1[6]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[24] <= ((((((main_crc32_inserter_last[16] ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[25] <= ((((main_crc32_inserter_last[17] ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]);
	main_crc32_inserter_next[26] <= ((((((((main_crc32_inserter_last[18] ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]) ^ main_crc32_inserter_last[24]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_data1[7]);
	main_crc32_inserter_next[27] <= ((((((((main_crc32_inserter_last[19] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]) ^ main_crc32_inserter_last[25]) ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_data1[6]);
	main_crc32_inserter_next[28] <= ((((((main_crc32_inserter_last[20] ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]) ^ main_crc32_inserter_last[26]) ^ main_crc32_inserter_data1[5]);
	main_crc32_inserter_next[29] <= ((((((main_crc32_inserter_last[21] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[30]) ^ main_crc32_inserter_data1[1]) ^ main_crc32_inserter_last[27]) ^ main_crc32_inserter_data1[4]);
	main_crc32_inserter_next[30] <= ((((main_crc32_inserter_last[22] ^ main_crc32_inserter_last[31]) ^ main_crc32_inserter_data1[0]) ^ main_crc32_inserter_last[28]) ^ main_crc32_inserter_data1[3]);
	main_crc32_inserter_next[31] <= ((main_crc32_inserter_last[23] ^ main_crc32_inserter_last[29]) ^ main_crc32_inserter_data1[2]);
// synthesis translate_off
	dummy_d_33 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_34;
// synthesis translate_on
always @(*) begin
	main_crc32_inserter_sink_ack <= 1'd0;
	main_crc32_inserter_source_stb <= 1'd0;
	main_crc32_inserter_source_eop <= 1'd0;
	main_crc32_inserter_source_payload_data <= 8'd0;
	main_crc32_inserter_source_payload_last_be <= 1'd0;
	main_crc32_inserter_source_payload_error <= 1'd0;
	main_crc32_inserter_data0 <= 8'd0;
	main_crc32_inserter_ce <= 1'd0;
	main_crc32_inserter_reset <= 1'd0;
	main_crc32_inserter_is_ongoing0 <= 1'd0;
	main_crc32_inserter_is_ongoing1 <= 1'd0;
	builder_liteethmaccrc32inserter_next_state <= 2'd0;
	builder_liteethmaccrc32inserter_next_state <= builder_liteethmaccrc32inserter_state;
	case (builder_liteethmaccrc32inserter_state)
		1'd1: begin
			main_crc32_inserter_ce <= (main_crc32_inserter_sink_stb & main_crc32_inserter_source_ack);
			main_crc32_inserter_data0 <= main_crc32_inserter_sink_payload_data;
			main_crc32_inserter_source_stb <= main_crc32_inserter_sink_stb;
			main_crc32_inserter_sink_ack <= main_crc32_inserter_source_ack;
			main_crc32_inserter_source_eop <= main_crc32_inserter_sink_eop;
			main_crc32_inserter_source_payload_data <= main_crc32_inserter_sink_payload_data;
			main_crc32_inserter_source_payload_last_be <= main_crc32_inserter_sink_payload_last_be;
			main_crc32_inserter_source_payload_error <= main_crc32_inserter_sink_payload_error;
			main_crc32_inserter_source_eop <= 1'd0;
			if (((main_crc32_inserter_sink_stb & main_crc32_inserter_sink_eop) & main_crc32_inserter_source_ack)) begin
				builder_liteethmaccrc32inserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_crc32_inserter_source_stb <= 1'd1;
			case (main_crc32_inserter_cnt)
				1'd0: begin
					main_crc32_inserter_source_payload_data <= main_crc32_inserter_value[31:24];
				end
				1'd1: begin
					main_crc32_inserter_source_payload_data <= main_crc32_inserter_value[23:16];
				end
				2'd2: begin
					main_crc32_inserter_source_payload_data <= main_crc32_inserter_value[15:8];
				end
				default: begin
					main_crc32_inserter_source_payload_data <= main_crc32_inserter_value[7:0];
				end
			endcase
			if (main_crc32_inserter_cnt_done) begin
				main_crc32_inserter_source_eop <= 1'd1;
				if (main_crc32_inserter_source_ack) begin
					builder_liteethmaccrc32inserter_next_state <= 1'd0;
				end
			end
			main_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			main_crc32_inserter_reset <= 1'd1;
			main_crc32_inserter_sink_ack <= 1'd1;
			if (main_crc32_inserter_sink_stb) begin
				main_crc32_inserter_sink_ack <= 1'd0;
				builder_liteethmaccrc32inserter_next_state <= 1'd1;
			end
			main_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_34 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_checker_fifo_full = (main_crc32_checker_syncfifo_level == 3'd4);
assign main_crc32_checker_fifo_in = (main_crc32_checker_sink_sink_stb & ((~main_crc32_checker_fifo_full) | main_crc32_checker_fifo_out));
assign main_crc32_checker_fifo_out = (main_crc32_checker_source_source_stb & main_crc32_checker_source_source_ack);
assign main_crc32_checker_syncfifo_sink_eop = main_crc32_checker_sink_sink_eop;
assign main_crc32_checker_syncfifo_sink_payload_data = main_crc32_checker_sink_sink_payload_data;
assign main_crc32_checker_syncfifo_sink_payload_last_be = main_crc32_checker_sink_sink_payload_last_be;
assign main_crc32_checker_syncfifo_sink_payload_error = main_crc32_checker_sink_sink_payload_error;

// synthesis translate_off
reg dummy_d_35;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_syncfifo_sink_stb <= 1'd0;
	main_crc32_checker_syncfifo_sink_stb <= main_crc32_checker_sink_sink_stb;
	main_crc32_checker_syncfifo_sink_stb <= main_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_35 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_36;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_sink_sink_ack <= 1'd0;
	main_crc32_checker_sink_sink_ack <= main_crc32_checker_syncfifo_sink_ack;
	main_crc32_checker_sink_sink_ack <= main_crc32_checker_fifo_in;
// synthesis translate_off
	dummy_d_36 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_checker_source_source_stb = (main_crc32_checker_sink_sink_stb & main_crc32_checker_fifo_full);
assign main_crc32_checker_source_source_eop = main_crc32_checker_sink_sink_eop;
assign main_crc32_checker_syncfifo_source_ack = main_crc32_checker_fifo_out;
assign main_crc32_checker_source_source_payload_data = main_crc32_checker_syncfifo_source_payload_data;
assign main_crc32_checker_source_source_payload_last_be = main_crc32_checker_syncfifo_source_payload_last_be;

// synthesis translate_off
reg dummy_d_37;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_source_source_payload_error <= 1'd0;
	main_crc32_checker_source_source_payload_error <= main_crc32_checker_syncfifo_source_payload_error;
	main_crc32_checker_source_source_payload_error <= (main_crc32_checker_sink_sink_payload_error | main_crc32_checker_crc_error);
// synthesis translate_off
	dummy_d_37 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_checker_error = ((main_crc32_checker_source_source_stb & main_crc32_checker_source_source_eop) & main_crc32_checker_crc_error);
assign main_crc32_checker_crc_data0 = main_crc32_checker_sink_sink_payload_data;
assign main_crc32_checker_crc_data1 = main_crc32_checker_crc_data0;
assign main_crc32_checker_crc_last = main_crc32_checker_crc_reg;
assign main_crc32_checker_crc_value = (~{main_crc32_checker_crc_reg[0], main_crc32_checker_crc_reg[1], main_crc32_checker_crc_reg[2], main_crc32_checker_crc_reg[3], main_crc32_checker_crc_reg[4], main_crc32_checker_crc_reg[5], main_crc32_checker_crc_reg[6], main_crc32_checker_crc_reg[7], main_crc32_checker_crc_reg[8], main_crc32_checker_crc_reg[9], main_crc32_checker_crc_reg[10], main_crc32_checker_crc_reg[11], main_crc32_checker_crc_reg[12], main_crc32_checker_crc_reg[13], main_crc32_checker_crc_reg[14], main_crc32_checker_crc_reg[15], main_crc32_checker_crc_reg[16], main_crc32_checker_crc_reg[17], main_crc32_checker_crc_reg[18], main_crc32_checker_crc_reg[19], main_crc32_checker_crc_reg[20], main_crc32_checker_crc_reg[21], main_crc32_checker_crc_reg[22], main_crc32_checker_crc_reg[23], main_crc32_checker_crc_reg[24], main_crc32_checker_crc_reg[25], main_crc32_checker_crc_reg[26], main_crc32_checker_crc_reg[27], main_crc32_checker_crc_reg[28], main_crc32_checker_crc_reg[29], main_crc32_checker_crc_reg[30], main_crc32_checker_crc_reg[31]});
assign main_crc32_checker_crc_error = (main_crc32_checker_crc_next != 32'd3338984827);

// synthesis translate_off
reg dummy_d_38;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_crc_next <= 32'd0;
	main_crc32_checker_crc_next[0] <= (((main_crc32_checker_crc_last[24] ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[1] <= (((((((main_crc32_checker_crc_last[25] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[2] <= (((((((((main_crc32_checker_crc_last[26] ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[3] <= (((((((main_crc32_checker_crc_last[27] ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[4] <= (((((((((main_crc32_checker_crc_last[28] ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[5] <= (((((((((((((main_crc32_checker_crc_last[29] ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[6] <= (((((((((((main_crc32_checker_crc_last[30] ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[7] <= (((((((((main_crc32_checker_crc_last[31] ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[8] <= ((((((((main_crc32_checker_crc_last[0] ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[9] <= ((((((((main_crc32_checker_crc_last[1] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[10] <= ((((((((main_crc32_checker_crc_last[2] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[11] <= ((((((((main_crc32_checker_crc_last[3] ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[12] <= ((((((((((((main_crc32_checker_crc_last[4] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[13] <= ((((((((((((main_crc32_checker_crc_last[5] ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[14] <= ((((((((((main_crc32_checker_crc_last[6] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]);
	main_crc32_checker_crc_next[15] <= ((((((((main_crc32_checker_crc_last[7] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]);
	main_crc32_checker_crc_next[16] <= ((((((main_crc32_checker_crc_last[8] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[17] <= ((((((main_crc32_checker_crc_last[9] ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[18] <= ((((((main_crc32_checker_crc_last[10] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]);
	main_crc32_checker_crc_next[19] <= ((((main_crc32_checker_crc_last[11] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]);
	main_crc32_checker_crc_next[20] <= ((main_crc32_checker_crc_last[12] ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]);
	main_crc32_checker_crc_next[21] <= ((main_crc32_checker_crc_last[13] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]);
	main_crc32_checker_crc_next[22] <= ((main_crc32_checker_crc_last[14] ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[23] <= ((((((main_crc32_checker_crc_last[15] ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_data1[6]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[24] <= ((((((main_crc32_checker_crc_last[16] ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[25] <= ((((main_crc32_checker_crc_last[17] ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]);
	main_crc32_checker_crc_next[26] <= ((((((((main_crc32_checker_crc_last[18] ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]) ^ main_crc32_checker_crc_last[24]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_data1[7]);
	main_crc32_checker_crc_next[27] <= ((((((((main_crc32_checker_crc_last[19] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]) ^ main_crc32_checker_crc_last[25]) ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_data1[6]);
	main_crc32_checker_crc_next[28] <= ((((((main_crc32_checker_crc_last[20] ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]) ^ main_crc32_checker_crc_last[26]) ^ main_crc32_checker_crc_data1[5]);
	main_crc32_checker_crc_next[29] <= ((((((main_crc32_checker_crc_last[21] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[30]) ^ main_crc32_checker_crc_data1[1]) ^ main_crc32_checker_crc_last[27]) ^ main_crc32_checker_crc_data1[4]);
	main_crc32_checker_crc_next[30] <= ((((main_crc32_checker_crc_last[22] ^ main_crc32_checker_crc_last[31]) ^ main_crc32_checker_crc_data1[0]) ^ main_crc32_checker_crc_last[28]) ^ main_crc32_checker_crc_data1[3]);
	main_crc32_checker_crc_next[31] <= ((main_crc32_checker_crc_last[23] ^ main_crc32_checker_crc_last[29]) ^ main_crc32_checker_crc_data1[2]);
// synthesis translate_off
	dummy_d_38 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_checker_syncfifo_syncfifo_din = {main_crc32_checker_syncfifo_fifo_in_eop, main_crc32_checker_syncfifo_fifo_in_payload_error, main_crc32_checker_syncfifo_fifo_in_payload_last_be, main_crc32_checker_syncfifo_fifo_in_payload_data};
assign {main_crc32_checker_syncfifo_fifo_out_eop, main_crc32_checker_syncfifo_fifo_out_payload_error, main_crc32_checker_syncfifo_fifo_out_payload_last_be, main_crc32_checker_syncfifo_fifo_out_payload_data} = main_crc32_checker_syncfifo_syncfifo_dout;
assign main_crc32_checker_syncfifo_sink_ack = main_crc32_checker_syncfifo_syncfifo_writable;
assign main_crc32_checker_syncfifo_syncfifo_we = main_crc32_checker_syncfifo_sink_stb;
assign main_crc32_checker_syncfifo_fifo_in_eop = main_crc32_checker_syncfifo_sink_eop;
assign main_crc32_checker_syncfifo_fifo_in_payload_data = main_crc32_checker_syncfifo_sink_payload_data;
assign main_crc32_checker_syncfifo_fifo_in_payload_last_be = main_crc32_checker_syncfifo_sink_payload_last_be;
assign main_crc32_checker_syncfifo_fifo_in_payload_error = main_crc32_checker_syncfifo_sink_payload_error;
assign main_crc32_checker_syncfifo_source_stb = main_crc32_checker_syncfifo_syncfifo_readable;
assign main_crc32_checker_syncfifo_source_eop = main_crc32_checker_syncfifo_fifo_out_eop;
assign main_crc32_checker_syncfifo_source_payload_data = main_crc32_checker_syncfifo_fifo_out_payload_data;
assign main_crc32_checker_syncfifo_source_payload_last_be = main_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign main_crc32_checker_syncfifo_source_payload_error = main_crc32_checker_syncfifo_fifo_out_payload_error;
assign main_crc32_checker_syncfifo_syncfifo_re = main_crc32_checker_syncfifo_source_ack;

// synthesis translate_off
reg dummy_d_39;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (main_crc32_checker_syncfifo_replace) begin
		main_crc32_checker_syncfifo_wrport_adr <= (main_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		main_crc32_checker_syncfifo_wrport_adr <= main_crc32_checker_syncfifo_produce;
	end
// synthesis translate_off
	dummy_d_39 <= dummy_s;
// synthesis translate_on
end
assign main_crc32_checker_syncfifo_wrport_dat_w = main_crc32_checker_syncfifo_syncfifo_din;
assign main_crc32_checker_syncfifo_wrport_we = (main_crc32_checker_syncfifo_syncfifo_we & (main_crc32_checker_syncfifo_syncfifo_writable | main_crc32_checker_syncfifo_replace));
assign main_crc32_checker_syncfifo_do_read = (main_crc32_checker_syncfifo_syncfifo_readable & main_crc32_checker_syncfifo_syncfifo_re);
assign main_crc32_checker_syncfifo_rdport_adr = main_crc32_checker_syncfifo_consume;
assign main_crc32_checker_syncfifo_syncfifo_dout = main_crc32_checker_syncfifo_rdport_dat_r;
assign main_crc32_checker_syncfifo_syncfifo_writable = (main_crc32_checker_syncfifo_level != 3'd5);
assign main_crc32_checker_syncfifo_syncfifo_readable = (main_crc32_checker_syncfifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_40;
// synthesis translate_on
always @(*) begin
	main_crc32_checker_crc_ce <= 1'd0;
	main_crc32_checker_crc_reset <= 1'd0;
	main_crc32_checker_fifo_reset <= 1'd0;
	builder_liteethmaccrc32checker_next_state <= 2'd0;
	builder_liteethmaccrc32checker_next_state <= builder_liteethmaccrc32checker_state;
	case (builder_liteethmaccrc32checker_state)
		1'd1: begin
			if ((main_crc32_checker_sink_sink_stb & main_crc32_checker_sink_sink_ack)) begin
				main_crc32_checker_crc_ce <= 1'd1;
				builder_liteethmaccrc32checker_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((main_crc32_checker_sink_sink_stb & main_crc32_checker_sink_sink_ack)) begin
				main_crc32_checker_crc_ce <= 1'd1;
				if (main_crc32_checker_sink_sink_eop) begin
					builder_liteethmaccrc32checker_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_crc32_checker_crc_reset <= 1'd1;
			main_crc32_checker_fifo_reset <= 1'd1;
			builder_liteethmaccrc32checker_next_state <= 1'd1;
		end
	endcase
// synthesis translate_off
	dummy_d_40 <= dummy_s;
// synthesis translate_on
end
assign main_ps_preamble_error_o = (main_ps_preamble_error_toggle_o ^ main_ps_preamble_error_toggle_o_r);
assign main_ps_crc_error_o = (main_ps_crc_error_toggle_o ^ main_ps_crc_error_toggle_o_r);
assign main_padding_inserter_counter_done = (main_padding_inserter_counter >= 6'd59);

// synthesis translate_off
reg dummy_d_41;
// synthesis translate_on
always @(*) begin
	main_padding_inserter_sink_ack <= 1'd0;
	main_padding_inserter_source_stb <= 1'd0;
	main_padding_inserter_source_eop <= 1'd0;
	main_padding_inserter_source_payload_data <= 8'd0;
	main_padding_inserter_source_payload_last_be <= 1'd0;
	main_padding_inserter_source_payload_error <= 1'd0;
	main_padding_inserter_counter_reset <= 1'd0;
	main_padding_inserter_counter_ce <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= 1'd0;
	builder_liteethmacpaddinginserter_next_state <= builder_liteethmacpaddinginserter_state;
	case (builder_liteethmacpaddinginserter_state)
		1'd1: begin
			main_padding_inserter_source_stb <= 1'd1;
			main_padding_inserter_source_eop <= main_padding_inserter_counter_done;
			main_padding_inserter_source_payload_data <= 1'd0;
			if ((main_padding_inserter_source_stb & main_padding_inserter_source_ack)) begin
				main_padding_inserter_counter_ce <= 1'd1;
				if (main_padding_inserter_counter_done) begin
					main_padding_inserter_counter_reset <= 1'd1;
					builder_liteethmacpaddinginserter_next_state <= 1'd0;
				end
			end
		end
		default: begin
			main_padding_inserter_source_stb <= main_padding_inserter_sink_stb;
			main_padding_inserter_sink_ack <= main_padding_inserter_source_ack;
			main_padding_inserter_source_eop <= main_padding_inserter_sink_eop;
			main_padding_inserter_source_payload_data <= main_padding_inserter_sink_payload_data;
			main_padding_inserter_source_payload_last_be <= main_padding_inserter_sink_payload_last_be;
			main_padding_inserter_source_payload_error <= main_padding_inserter_sink_payload_error;
			if ((main_padding_inserter_source_stb & main_padding_inserter_source_ack)) begin
				main_padding_inserter_counter_ce <= 1'd1;
				if (main_padding_inserter_sink_eop) begin
					if ((~main_padding_inserter_counter_done)) begin
						main_padding_inserter_source_eop <= 1'd0;
						builder_liteethmacpaddinginserter_next_state <= 1'd1;
					end else begin
						main_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_41 <= dummy_s;
// synthesis translate_on
end
assign main_padding_checker_source_stb = main_padding_checker_sink_stb;
assign main_padding_checker_sink_ack = main_padding_checker_source_ack;
assign main_padding_checker_source_eop = main_padding_checker_sink_eop;
assign main_padding_checker_source_payload_data = main_padding_checker_sink_payload_data;
assign main_padding_checker_source_payload_last_be = main_padding_checker_sink_payload_last_be;
assign main_padding_checker_source_payload_error = main_padding_checker_sink_payload_error;
assign main_tx_last_be_source_stb = (main_tx_last_be_sink_stb & main_tx_last_be_ongoing);
assign main_tx_last_be_source_eop = main_tx_last_be_sink_payload_last_be;
assign main_tx_last_be_source_payload_data = main_tx_last_be_sink_payload_data;
assign main_tx_last_be_sink_ack = main_tx_last_be_source_ack;
assign main_rx_last_be_source_stb = main_rx_last_be_sink_stb;
assign main_rx_last_be_sink_ack = main_rx_last_be_source_ack;
assign main_rx_last_be_source_eop = main_rx_last_be_sink_eop;
assign main_rx_last_be_source_payload_data = main_rx_last_be_sink_payload_data;
assign main_rx_last_be_source_payload_error = main_rx_last_be_sink_payload_error;

// synthesis translate_off
reg dummy_d_42;
// synthesis translate_on
always @(*) begin
	main_rx_last_be_source_payload_last_be <= 1'd0;
	main_rx_last_be_source_payload_last_be <= main_rx_last_be_sink_payload_last_be;
	main_rx_last_be_source_payload_last_be <= main_rx_last_be_sink_eop;
// synthesis translate_off
	dummy_d_42 <= dummy_s;
// synthesis translate_on
end
assign main_tx_converter_converter_sink_stb = main_tx_converter_sink_sink_stb;
assign main_tx_converter_converter_sink_eop = main_tx_converter_sink_sink_eop;
assign main_tx_converter_sink_sink_ack = main_tx_converter_converter_sink_ack;

// synthesis translate_off
reg dummy_d_43;
// synthesis translate_on
always @(*) begin
	main_tx_converter_converter_sink_payload_data <= 40'd0;
	main_tx_converter_converter_sink_payload_data[7:0] <= main_tx_converter_sink_sink_payload_data[7:0];
	main_tx_converter_converter_sink_payload_data[8] <= main_tx_converter_sink_sink_payload_last_be[0];
	main_tx_converter_converter_sink_payload_data[9] <= main_tx_converter_sink_sink_payload_error[0];
	main_tx_converter_converter_sink_payload_data[17:10] <= main_tx_converter_sink_sink_payload_data[15:8];
	main_tx_converter_converter_sink_payload_data[18] <= main_tx_converter_sink_sink_payload_last_be[1];
	main_tx_converter_converter_sink_payload_data[19] <= main_tx_converter_sink_sink_payload_error[1];
	main_tx_converter_converter_sink_payload_data[27:20] <= main_tx_converter_sink_sink_payload_data[23:16];
	main_tx_converter_converter_sink_payload_data[28] <= main_tx_converter_sink_sink_payload_last_be[2];
	main_tx_converter_converter_sink_payload_data[29] <= main_tx_converter_sink_sink_payload_error[2];
	main_tx_converter_converter_sink_payload_data[37:30] <= main_tx_converter_sink_sink_payload_data[31:24];
	main_tx_converter_converter_sink_payload_data[38] <= main_tx_converter_sink_sink_payload_last_be[3];
	main_tx_converter_converter_sink_payload_data[39] <= main_tx_converter_sink_sink_payload_error[3];
// synthesis translate_off
	dummy_d_43 <= dummy_s;
// synthesis translate_on
end
assign main_tx_converter_source_source_stb = main_tx_converter_converter_source_stb;
assign main_tx_converter_source_source_eop = main_tx_converter_converter_source_eop;
assign main_tx_converter_converter_source_ack = main_tx_converter_source_source_ack;
assign {main_tx_converter_source_source_payload_error, main_tx_converter_source_source_payload_last_be, main_tx_converter_source_source_payload_data} = main_tx_converter_converter_source_payload_data;
assign main_tx_converter_converter_last = (main_tx_converter_converter_mux == 2'd3);
assign main_tx_converter_converter_source_stb = main_tx_converter_converter_sink_stb;
assign main_tx_converter_converter_source_eop = (main_tx_converter_converter_sink_eop & main_tx_converter_converter_last);
assign main_tx_converter_converter_sink_ack = (main_tx_converter_converter_last & main_tx_converter_converter_source_ack);

// synthesis translate_off
reg dummy_d_44;
// synthesis translate_on
always @(*) begin
	main_tx_converter_converter_source_payload_data <= 10'd0;
	case (main_tx_converter_converter_mux)
		1'd0: begin
			main_tx_converter_converter_source_payload_data <= main_tx_converter_converter_sink_payload_data[39:30];
		end
		1'd1: begin
			main_tx_converter_converter_source_payload_data <= main_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd2: begin
			main_tx_converter_converter_source_payload_data <= main_tx_converter_converter_sink_payload_data[19:10];
		end
		default: begin
			main_tx_converter_converter_source_payload_data <= main_tx_converter_converter_sink_payload_data[9:0];
		end
	endcase
// synthesis translate_off
	dummy_d_44 <= dummy_s;
// synthesis translate_on
end
assign main_rx_converter_converter_sink_stb = main_rx_converter_sink_sink_stb;
assign main_rx_converter_converter_sink_eop = main_rx_converter_sink_sink_eop;
assign main_rx_converter_sink_sink_ack = main_rx_converter_converter_sink_ack;
assign main_rx_converter_converter_sink_payload_data = {main_rx_converter_sink_sink_payload_error, main_rx_converter_sink_sink_payload_last_be, main_rx_converter_sink_sink_payload_data};
assign main_rx_converter_source_source_stb = main_rx_converter_converter_source_stb;
assign main_rx_converter_source_source_eop = main_rx_converter_converter_source_eop;
assign main_rx_converter_converter_source_ack = main_rx_converter_source_source_ack;

// synthesis translate_off
reg dummy_d_45;
// synthesis translate_on
always @(*) begin
	main_rx_converter_source_source_payload_data <= 32'd0;
	main_rx_converter_source_source_payload_data[7:0] <= main_rx_converter_converter_source_payload_data[7:0];
	main_rx_converter_source_source_payload_data[15:8] <= main_rx_converter_converter_source_payload_data[17:10];
	main_rx_converter_source_source_payload_data[23:16] <= main_rx_converter_converter_source_payload_data[27:20];
	main_rx_converter_source_source_payload_data[31:24] <= main_rx_converter_converter_source_payload_data[37:30];
// synthesis translate_off
	dummy_d_45 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_46;
// synthesis translate_on
always @(*) begin
	main_rx_converter_source_source_payload_last_be <= 4'd0;
	main_rx_converter_source_source_payload_last_be[0] <= main_rx_converter_converter_source_payload_data[8];
	main_rx_converter_source_source_payload_last_be[1] <= main_rx_converter_converter_source_payload_data[18];
	main_rx_converter_source_source_payload_last_be[2] <= main_rx_converter_converter_source_payload_data[28];
	main_rx_converter_source_source_payload_last_be[3] <= main_rx_converter_converter_source_payload_data[38];
// synthesis translate_off
	dummy_d_46 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_47;
// synthesis translate_on
always @(*) begin
	main_rx_converter_source_source_payload_error <= 4'd0;
	main_rx_converter_source_source_payload_error[0] <= main_rx_converter_converter_source_payload_data[9];
	main_rx_converter_source_source_payload_error[1] <= main_rx_converter_converter_source_payload_data[19];
	main_rx_converter_source_source_payload_error[2] <= main_rx_converter_converter_source_payload_data[29];
	main_rx_converter_source_source_payload_error[3] <= main_rx_converter_converter_source_payload_data[39];
// synthesis translate_off
	dummy_d_47 <= dummy_s;
// synthesis translate_on
end
assign main_rx_converter_converter_sink_ack = ((~main_rx_converter_converter_strobe_all) | main_rx_converter_converter_source_ack);
assign main_rx_converter_converter_source_stb = main_rx_converter_converter_strobe_all;
assign main_rx_converter_converter_load_part = (main_rx_converter_converter_sink_stb & main_rx_converter_converter_sink_ack);
assign main_tx_cdc_asyncfifo_din = {main_tx_cdc_fifo_in_eop, main_tx_cdc_fifo_in_payload_error, main_tx_cdc_fifo_in_payload_last_be, main_tx_cdc_fifo_in_payload_data};
assign {main_tx_cdc_fifo_out_eop, main_tx_cdc_fifo_out_payload_error, main_tx_cdc_fifo_out_payload_last_be, main_tx_cdc_fifo_out_payload_data} = main_tx_cdc_asyncfifo_dout;
assign main_tx_cdc_sink_ack = main_tx_cdc_asyncfifo_writable;
assign main_tx_cdc_asyncfifo_we = main_tx_cdc_sink_stb;
assign main_tx_cdc_fifo_in_eop = main_tx_cdc_sink_eop;
assign main_tx_cdc_fifo_in_payload_data = main_tx_cdc_sink_payload_data;
assign main_tx_cdc_fifo_in_payload_last_be = main_tx_cdc_sink_payload_last_be;
assign main_tx_cdc_fifo_in_payload_error = main_tx_cdc_sink_payload_error;
assign main_tx_cdc_source_stb = main_tx_cdc_asyncfifo_readable;
assign main_tx_cdc_source_eop = main_tx_cdc_fifo_out_eop;
assign main_tx_cdc_source_payload_data = main_tx_cdc_fifo_out_payload_data;
assign main_tx_cdc_source_payload_last_be = main_tx_cdc_fifo_out_payload_last_be;
assign main_tx_cdc_source_payload_error = main_tx_cdc_fifo_out_payload_error;
assign main_tx_cdc_asyncfifo_re = main_tx_cdc_source_ack;
assign main_tx_cdc_graycounter0_ce = (main_tx_cdc_asyncfifo_writable & main_tx_cdc_asyncfifo_we);
assign main_tx_cdc_graycounter1_ce = (main_tx_cdc_asyncfifo_readable & main_tx_cdc_asyncfifo_re);
assign main_tx_cdc_asyncfifo_writable = (((main_tx_cdc_graycounter0_q[6] == main_tx_cdc_consume_wdomain[6]) | (main_tx_cdc_graycounter0_q[5] == main_tx_cdc_consume_wdomain[5])) | (main_tx_cdc_graycounter0_q[4:0] != main_tx_cdc_consume_wdomain[4:0]));
assign main_tx_cdc_asyncfifo_readable = (main_tx_cdc_graycounter1_q != main_tx_cdc_produce_rdomain);
assign main_tx_cdc_wrport_adr = main_tx_cdc_graycounter0_q_binary[5:0];
assign main_tx_cdc_wrport_dat_w = main_tx_cdc_asyncfifo_din;
assign main_tx_cdc_wrport_we = main_tx_cdc_graycounter0_ce;
assign main_tx_cdc_rdport_adr = main_tx_cdc_graycounter1_q_next_binary[5:0];
assign main_tx_cdc_asyncfifo_dout = main_tx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_48;
// synthesis translate_on
always @(*) begin
	main_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_tx_cdc_graycounter0_ce) begin
		main_tx_cdc_graycounter0_q_next_binary <= (main_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_tx_cdc_graycounter0_q_next_binary <= main_tx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_48 <= dummy_s;
// synthesis translate_on
end
assign main_tx_cdc_graycounter0_q_next = (main_tx_cdc_graycounter0_q_next_binary ^ main_tx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_49;
// synthesis translate_on
always @(*) begin
	main_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_tx_cdc_graycounter1_ce) begin
		main_tx_cdc_graycounter1_q_next_binary <= (main_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_tx_cdc_graycounter1_q_next_binary <= main_tx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_49 <= dummy_s;
// synthesis translate_on
end
assign main_tx_cdc_graycounter1_q_next = (main_tx_cdc_graycounter1_q_next_binary ^ main_tx_cdc_graycounter1_q_next_binary[6:1]);
assign main_rx_cdc_asyncfifo_din = {main_rx_cdc_fifo_in_eop, main_rx_cdc_fifo_in_payload_error, main_rx_cdc_fifo_in_payload_last_be, main_rx_cdc_fifo_in_payload_data};
assign {main_rx_cdc_fifo_out_eop, main_rx_cdc_fifo_out_payload_error, main_rx_cdc_fifo_out_payload_last_be, main_rx_cdc_fifo_out_payload_data} = main_rx_cdc_asyncfifo_dout;
assign main_rx_cdc_sink_ack = main_rx_cdc_asyncfifo_writable;
assign main_rx_cdc_asyncfifo_we = main_rx_cdc_sink_stb;
assign main_rx_cdc_fifo_in_eop = main_rx_cdc_sink_eop;
assign main_rx_cdc_fifo_in_payload_data = main_rx_cdc_sink_payload_data;
assign main_rx_cdc_fifo_in_payload_last_be = main_rx_cdc_sink_payload_last_be;
assign main_rx_cdc_fifo_in_payload_error = main_rx_cdc_sink_payload_error;
assign main_rx_cdc_source_stb = main_rx_cdc_asyncfifo_readable;
assign main_rx_cdc_source_eop = main_rx_cdc_fifo_out_eop;
assign main_rx_cdc_source_payload_data = main_rx_cdc_fifo_out_payload_data;
assign main_rx_cdc_source_payload_last_be = main_rx_cdc_fifo_out_payload_last_be;
assign main_rx_cdc_source_payload_error = main_rx_cdc_fifo_out_payload_error;
assign main_rx_cdc_asyncfifo_re = main_rx_cdc_source_ack;
assign main_rx_cdc_graycounter0_ce = (main_rx_cdc_asyncfifo_writable & main_rx_cdc_asyncfifo_we);
assign main_rx_cdc_graycounter1_ce = (main_rx_cdc_asyncfifo_readable & main_rx_cdc_asyncfifo_re);
assign main_rx_cdc_asyncfifo_writable = (((main_rx_cdc_graycounter0_q[6] == main_rx_cdc_consume_wdomain[6]) | (main_rx_cdc_graycounter0_q[5] == main_rx_cdc_consume_wdomain[5])) | (main_rx_cdc_graycounter0_q[4:0] != main_rx_cdc_consume_wdomain[4:0]));
assign main_rx_cdc_asyncfifo_readable = (main_rx_cdc_graycounter1_q != main_rx_cdc_produce_rdomain);
assign main_rx_cdc_wrport_adr = main_rx_cdc_graycounter0_q_binary[5:0];
assign main_rx_cdc_wrport_dat_w = main_rx_cdc_asyncfifo_din;
assign main_rx_cdc_wrport_we = main_rx_cdc_graycounter0_ce;
assign main_rx_cdc_rdport_adr = main_rx_cdc_graycounter1_q_next_binary[5:0];
assign main_rx_cdc_asyncfifo_dout = main_rx_cdc_rdport_dat_r;

// synthesis translate_off
reg dummy_d_50;
// synthesis translate_on
always @(*) begin
	main_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (main_rx_cdc_graycounter0_ce) begin
		main_rx_cdc_graycounter0_q_next_binary <= (main_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		main_rx_cdc_graycounter0_q_next_binary <= main_rx_cdc_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_50 <= dummy_s;
// synthesis translate_on
end
assign main_rx_cdc_graycounter0_q_next = (main_rx_cdc_graycounter0_q_next_binary ^ main_rx_cdc_graycounter0_q_next_binary[6:1]);

// synthesis translate_off
reg dummy_d_51;
// synthesis translate_on
always @(*) begin
	main_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (main_rx_cdc_graycounter1_ce) begin
		main_rx_cdc_graycounter1_q_next_binary <= (main_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		main_rx_cdc_graycounter1_q_next_binary <= main_rx_cdc_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_51 <= dummy_s;
// synthesis translate_on
end
assign main_rx_cdc_graycounter1_q_next = (main_rx_cdc_graycounter1_q_next_binary ^ main_rx_cdc_graycounter1_q_next_binary[6:1]);
assign main_writer_sink_sink_stb = main_sink_stb;
assign main_sink_ack = main_writer_sink_sink_ack;
assign main_writer_sink_sink_eop = main_sink_eop;
assign main_writer_sink_sink_payload_data = main_sink_payload_data;
assign main_writer_sink_sink_payload_last_be = main_sink_payload_last_be;
assign main_writer_sink_sink_payload_error = main_sink_payload_error;
assign main_source_stb = main_reader_source_source_stb;
assign main_reader_source_source_ack = main_source_ack;
assign main_source_eop = main_reader_source_source_eop;
assign main_source_payload_data = main_reader_source_source_payload_data;
assign main_source_payload_last_be = main_reader_source_source_payload_last_be;
assign main_source_payload_error = main_reader_source_source_payload_error;

// synthesis translate_off
reg dummy_d_52;
// synthesis translate_on
always @(*) begin
	main_writer_increment <= 3'd0;
	if (main_writer_sink_sink_payload_last_be[3]) begin
		main_writer_increment <= 1'd1;
	end else begin
		if (main_writer_sink_sink_payload_last_be[2]) begin
			main_writer_increment <= 2'd2;
		end else begin
			if (main_writer_sink_sink_payload_last_be[1]) begin
				main_writer_increment <= 2'd3;
			end else begin
				main_writer_increment <= 3'd4;
			end
		end
	end
// synthesis translate_off
	dummy_d_52 <= dummy_s;
// synthesis translate_on
end
assign main_writer_fifo_sink_payload_slot = main_writer_slot;
assign main_writer_fifo_sink_payload_length = main_writer_counter;
assign main_writer_fifo_source_ack = main_writer_available_clear;
assign main_writer_available_trigger = main_writer_fifo_source_stb;
assign main_writer_slot_status = main_writer_fifo_source_payload_slot;
assign main_writer_length_status = main_writer_fifo_source_payload_length;

// synthesis translate_off
reg dummy_d_53;
// synthesis translate_on
always @(*) begin
	main_writer_memory0_adr <= 9'd0;
	main_writer_memory0_we <= 1'd0;
	main_writer_memory0_dat_w <= 32'd0;
	main_writer_memory1_adr <= 9'd0;
	main_writer_memory1_we <= 1'd0;
	main_writer_memory1_dat_w <= 32'd0;
	main_writer_memory2_adr <= 9'd0;
	main_writer_memory2_we <= 1'd0;
	main_writer_memory2_dat_w <= 32'd0;
	main_writer_memory3_adr <= 9'd0;
	main_writer_memory3_we <= 1'd0;
	main_writer_memory3_dat_w <= 32'd0;
	case (main_writer_slot)
		1'd0: begin
			main_writer_memory0_adr <= main_writer_counter[31:2];
			main_writer_memory0_dat_w <= main_writer_sink_sink_payload_data;
			if ((main_writer_sink_sink_stb & main_writer_ongoing)) begin
				main_writer_memory0_we <= 4'd15;
			end
		end
		1'd1: begin
			main_writer_memory1_adr <= main_writer_counter[31:2];
			main_writer_memory1_dat_w <= main_writer_sink_sink_payload_data;
			if ((main_writer_sink_sink_stb & main_writer_ongoing)) begin
				main_writer_memory1_we <= 4'd15;
			end
		end
		2'd2: begin
			main_writer_memory2_adr <= main_writer_counter[31:2];
			main_writer_memory2_dat_w <= main_writer_sink_sink_payload_data;
			if ((main_writer_sink_sink_stb & main_writer_ongoing)) begin
				main_writer_memory2_we <= 4'd15;
			end
		end
		2'd3: begin
			main_writer_memory3_adr <= main_writer_counter[31:2];
			main_writer_memory3_dat_w <= main_writer_sink_sink_payload_data;
			if ((main_writer_sink_sink_stb & main_writer_ongoing)) begin
				main_writer_memory3_we <= 4'd15;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_53 <= dummy_s;
// synthesis translate_on
end
assign main_writer_status_w = main_writer_available_status;

// synthesis translate_off
reg dummy_d_54;
// synthesis translate_on
always @(*) begin
	main_writer_available_clear <= 1'd0;
	if ((main_writer_pending_re & main_writer_pending_r)) begin
		main_writer_available_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_54 <= dummy_s;
// synthesis translate_on
end
assign main_writer_pending_w = main_writer_available_pending;
assign main_writer_irq = (main_writer_pending_w & main_writer_storage);
assign main_writer_available_status = main_writer_available_trigger;
assign main_writer_available_pending = main_writer_available_trigger;
assign main_writer_fifo_syncfifo_din = {main_writer_fifo_fifo_in_eop, main_writer_fifo_fifo_in_payload_length, main_writer_fifo_fifo_in_payload_slot};
assign {main_writer_fifo_fifo_out_eop, main_writer_fifo_fifo_out_payload_length, main_writer_fifo_fifo_out_payload_slot} = main_writer_fifo_syncfifo_dout;
assign main_writer_fifo_sink_ack = main_writer_fifo_syncfifo_writable;
assign main_writer_fifo_syncfifo_we = main_writer_fifo_sink_stb;
assign main_writer_fifo_fifo_in_eop = main_writer_fifo_sink_eop;
assign main_writer_fifo_fifo_in_payload_slot = main_writer_fifo_sink_payload_slot;
assign main_writer_fifo_fifo_in_payload_length = main_writer_fifo_sink_payload_length;
assign main_writer_fifo_source_stb = main_writer_fifo_syncfifo_readable;
assign main_writer_fifo_source_eop = main_writer_fifo_fifo_out_eop;
assign main_writer_fifo_source_payload_slot = main_writer_fifo_fifo_out_payload_slot;
assign main_writer_fifo_source_payload_length = main_writer_fifo_fifo_out_payload_length;
assign main_writer_fifo_syncfifo_re = main_writer_fifo_source_ack;

// synthesis translate_off
reg dummy_d_55;
// synthesis translate_on
always @(*) begin
	main_writer_fifo_wrport_adr <= 2'd0;
	if (main_writer_fifo_replace) begin
		main_writer_fifo_wrport_adr <= (main_writer_fifo_produce - 1'd1);
	end else begin
		main_writer_fifo_wrport_adr <= main_writer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_55 <= dummy_s;
// synthesis translate_on
end
assign main_writer_fifo_wrport_dat_w = main_writer_fifo_syncfifo_din;
assign main_writer_fifo_wrport_we = (main_writer_fifo_syncfifo_we & (main_writer_fifo_syncfifo_writable | main_writer_fifo_replace));
assign main_writer_fifo_do_read = (main_writer_fifo_syncfifo_readable & main_writer_fifo_syncfifo_re);
assign main_writer_fifo_rdport_adr = main_writer_fifo_consume;
assign main_writer_fifo_syncfifo_dout = main_writer_fifo_rdport_dat_r;
assign main_writer_fifo_syncfifo_writable = (main_writer_fifo_level != 3'd4);
assign main_writer_fifo_syncfifo_readable = (main_writer_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_56;
// synthesis translate_on
always @(*) begin
	main_writer_counter_reset <= 1'd0;
	main_writer_counter_ce <= 1'd0;
	main_writer_slot_ce <= 1'd0;
	main_writer_ongoing <= 1'd0;
	main_writer_fifo_sink_stb <= 1'd0;
	builder_liteethmacsramwriter_next_state <= 2'd0;
	main_writer_errors_status_next_value <= 32'd0;
	main_writer_errors_status_next_value_ce <= 1'd0;
	builder_liteethmacsramwriter_next_state <= builder_liteethmacsramwriter_state;
	case (builder_liteethmacsramwriter_state)
		1'd1: begin
			if (main_writer_sink_sink_stb) begin
				if ((main_writer_counter == 11'd1530)) begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end else begin
					main_writer_counter_ce <= 1'd1;
					main_writer_ongoing <= 1'd1;
				end
				if (main_writer_sink_sink_eop) begin
					if (((main_writer_sink_sink_payload_error & main_writer_sink_sink_payload_last_be) != 1'd0)) begin
						main_writer_counter_reset <= 1'd1;
						builder_liteethmacsramwriter_next_state <= 1'd0;
					end else begin
						builder_liteethmacsramwriter_next_state <= 2'd3;
					end
				end
			end
		end
		2'd2: begin
			main_writer_counter_reset <= 1'd1;
			if ((main_writer_sink_sink_stb & main_writer_sink_sink_eop)) begin
				main_writer_errors_status_next_value <= (main_writer_errors_status + 1'd1);
				main_writer_errors_status_next_value_ce <= 1'd1;
				builder_liteethmacsramwriter_next_state <= 1'd0;
			end
		end
		2'd3: begin
			main_writer_counter_reset <= 1'd1;
			main_writer_slot_ce <= 1'd1;
			main_writer_fifo_sink_stb <= 1'd1;
			builder_liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (main_writer_sink_sink_stb) begin
				if (main_writer_fifo_sink_ack) begin
					main_writer_ongoing <= 1'd1;
					main_writer_counter_ce <= 1'd1;
					builder_liteethmacsramwriter_next_state <= 1'd1;
				end else begin
					builder_liteethmacsramwriter_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_56 <= dummy_s;
// synthesis translate_on
end
assign main_reader_fifo_sink_stb = main_reader_start_re;
assign main_reader_fifo_sink_payload_slot = main_reader_slot_storage;
assign main_reader_fifo_sink_payload_length = main_reader_length_storage;
assign main_reader_ready_status = main_reader_fifo_sink_ack;

// synthesis translate_off
reg dummy_d_57;
// synthesis translate_on
always @(*) begin
	main_reader_source_source_payload_last_be <= 4'd0;
	if (main_reader_last) begin
		if ((main_reader_fifo_source_payload_length[1:0] == 2'd3)) begin
			main_reader_source_source_payload_last_be <= 2'd2;
		end else begin
			if ((main_reader_fifo_source_payload_length[1:0] == 2'd2)) begin
				main_reader_source_source_payload_last_be <= 3'd4;
			end else begin
				if ((main_reader_fifo_source_payload_length[1:0] == 1'd1)) begin
					main_reader_source_source_payload_last_be <= 4'd8;
				end else begin
					main_reader_source_source_payload_last_be <= 1'd1;
				end
			end
		end
	end
// synthesis translate_off
	dummy_d_57 <= dummy_s;
// synthesis translate_on
end
assign main_reader_last = ((main_reader_counter + 3'd4) >= main_reader_fifo_source_payload_length);
assign main_reader_memory0_adr = main_reader_counter[10:2];
assign main_reader_memory1_adr = main_reader_counter[10:2];
assign main_reader_memory2_adr = main_reader_counter[10:2];
assign main_reader_memory3_adr = main_reader_counter[10:2];

// synthesis translate_off
reg dummy_d_58;
// synthesis translate_on
always @(*) begin
	main_reader_source_source_payload_data <= 32'd0;
	case (main_reader_fifo_source_payload_slot)
		1'd0: begin
			main_reader_source_source_payload_data <= main_reader_memory0_dat_r;
		end
		1'd1: begin
			main_reader_source_source_payload_data <= main_reader_memory1_dat_r;
		end
		2'd2: begin
			main_reader_source_source_payload_data <= main_reader_memory2_dat_r;
		end
		2'd3: begin
			main_reader_source_source_payload_data <= main_reader_memory3_dat_r;
		end
	endcase
// synthesis translate_off
	dummy_d_58 <= dummy_s;
// synthesis translate_on
end
assign main_reader_eventmanager_status_w = main_reader_done_status;

// synthesis translate_off
reg dummy_d_59;
// synthesis translate_on
always @(*) begin
	main_reader_done_clear <= 1'd0;
	if ((main_reader_eventmanager_pending_re & main_reader_eventmanager_pending_r)) begin
		main_reader_done_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_59 <= dummy_s;
// synthesis translate_on
end
assign main_reader_eventmanager_pending_w = main_reader_done_pending;
assign main_reader_irq = (main_reader_eventmanager_pending_w & main_reader_eventmanager_storage);
assign main_reader_done_status = 1'd0;
assign main_reader_fifo_syncfifo_din = {main_reader_fifo_fifo_in_eop, main_reader_fifo_fifo_in_payload_length, main_reader_fifo_fifo_in_payload_slot};
assign {main_reader_fifo_fifo_out_eop, main_reader_fifo_fifo_out_payload_length, main_reader_fifo_fifo_out_payload_slot} = main_reader_fifo_syncfifo_dout;
assign main_reader_fifo_sink_ack = main_reader_fifo_syncfifo_writable;
assign main_reader_fifo_syncfifo_we = main_reader_fifo_sink_stb;
assign main_reader_fifo_fifo_in_eop = main_reader_fifo_sink_eop;
assign main_reader_fifo_fifo_in_payload_slot = main_reader_fifo_sink_payload_slot;
assign main_reader_fifo_fifo_in_payload_length = main_reader_fifo_sink_payload_length;
assign main_reader_fifo_source_stb = main_reader_fifo_syncfifo_readable;
assign main_reader_fifo_source_eop = main_reader_fifo_fifo_out_eop;
assign main_reader_fifo_source_payload_slot = main_reader_fifo_fifo_out_payload_slot;
assign main_reader_fifo_source_payload_length = main_reader_fifo_fifo_out_payload_length;
assign main_reader_fifo_syncfifo_re = main_reader_fifo_source_ack;

// synthesis translate_off
reg dummy_d_60;
// synthesis translate_on
always @(*) begin
	main_reader_fifo_wrport_adr <= 2'd0;
	if (main_reader_fifo_replace) begin
		main_reader_fifo_wrport_adr <= (main_reader_fifo_produce - 1'd1);
	end else begin
		main_reader_fifo_wrport_adr <= main_reader_fifo_produce;
	end
// synthesis translate_off
	dummy_d_60 <= dummy_s;
// synthesis translate_on
end
assign main_reader_fifo_wrport_dat_w = main_reader_fifo_syncfifo_din;
assign main_reader_fifo_wrport_we = (main_reader_fifo_syncfifo_we & (main_reader_fifo_syncfifo_writable | main_reader_fifo_replace));
assign main_reader_fifo_do_read = (main_reader_fifo_syncfifo_readable & main_reader_fifo_syncfifo_re);
assign main_reader_fifo_rdport_adr = main_reader_fifo_consume;
assign main_reader_fifo_syncfifo_dout = main_reader_fifo_rdport_dat_r;
assign main_reader_fifo_syncfifo_writable = (main_reader_fifo_level != 3'd4);
assign main_reader_fifo_syncfifo_readable = (main_reader_fifo_level != 1'd0);

// synthesis translate_off
reg dummy_d_61;
// synthesis translate_on
always @(*) begin
	main_reader_source_source_stb <= 1'd0;
	main_reader_source_source_eop <= 1'd0;
	main_reader_done_trigger <= 1'd0;
	main_reader_fifo_source_ack <= 1'd0;
	main_reader_counter_reset <= 1'd0;
	main_reader_counter_ce <= 1'd0;
	builder_liteethmacsramreader_next_state <= 2'd0;
	builder_liteethmacsramreader_next_state <= builder_liteethmacsramreader_state;
	case (builder_liteethmacsramreader_state)
		1'd1: begin
			if ((~main_reader_last_d)) begin
				builder_liteethmacsramreader_next_state <= 2'd2;
			end else begin
				builder_liteethmacsramreader_next_state <= 2'd3;
			end
		end
		2'd2: begin
			main_reader_source_source_stb <= 1'd1;
			main_reader_source_source_eop <= main_reader_last;
			if (main_reader_source_source_ack) begin
				main_reader_counter_ce <= (~main_reader_last);
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
		2'd3: begin
			main_reader_fifo_source_ack <= 1'd1;
			main_reader_done_trigger <= 1'd1;
			builder_liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			main_reader_counter_reset <= 1'd1;
			if (main_reader_fifo_source_stb) begin
				builder_liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_61 <= dummy_s;
// synthesis translate_on
end
assign main_ev_irq = (main_writer_irq | main_reader_irq);
assign main_sram0_adr0 = main_sram0_bus_adr0[8:0];
assign main_sram0_bus_dat_r0 = main_sram0_dat_r0;
assign main_sram1_adr0 = main_sram1_bus_adr0[8:0];
assign main_sram1_bus_dat_r0 = main_sram1_dat_r0;
assign main_sram2_adr0 = main_sram2_bus_adr0[8:0];
assign main_sram2_bus_dat_r0 = main_sram2_dat_r0;
assign main_sram3_adr0 = main_sram3_bus_adr0[8:0];
assign main_sram3_bus_dat_r0 = main_sram3_dat_r0;

// synthesis translate_off
reg dummy_d_62;
// synthesis translate_on
always @(*) begin
	main_sram0_we <= 4'd0;
	main_sram0_we[0] <= (((main_sram0_bus_cyc1 & main_sram0_bus_stb1) & main_sram0_bus_we1) & main_sram0_bus_sel1[0]);
	main_sram0_we[1] <= (((main_sram0_bus_cyc1 & main_sram0_bus_stb1) & main_sram0_bus_we1) & main_sram0_bus_sel1[1]);
	main_sram0_we[2] <= (((main_sram0_bus_cyc1 & main_sram0_bus_stb1) & main_sram0_bus_we1) & main_sram0_bus_sel1[2]);
	main_sram0_we[3] <= (((main_sram0_bus_cyc1 & main_sram0_bus_stb1) & main_sram0_bus_we1) & main_sram0_bus_sel1[3]);
// synthesis translate_off
	dummy_d_62 <= dummy_s;
// synthesis translate_on
end
assign main_sram0_adr1 = main_sram0_bus_adr1[8:0];
assign main_sram0_bus_dat_r1 = main_sram0_dat_r1;
assign main_sram0_dat_w = main_sram0_bus_dat_w1;

// synthesis translate_off
reg dummy_d_63;
// synthesis translate_on
always @(*) begin
	main_sram1_we <= 4'd0;
	main_sram1_we[0] <= (((main_sram1_bus_cyc1 & main_sram1_bus_stb1) & main_sram1_bus_we1) & main_sram1_bus_sel1[0]);
	main_sram1_we[1] <= (((main_sram1_bus_cyc1 & main_sram1_bus_stb1) & main_sram1_bus_we1) & main_sram1_bus_sel1[1]);
	main_sram1_we[2] <= (((main_sram1_bus_cyc1 & main_sram1_bus_stb1) & main_sram1_bus_we1) & main_sram1_bus_sel1[2]);
	main_sram1_we[3] <= (((main_sram1_bus_cyc1 & main_sram1_bus_stb1) & main_sram1_bus_we1) & main_sram1_bus_sel1[3]);
// synthesis translate_off
	dummy_d_63 <= dummy_s;
// synthesis translate_on
end
assign main_sram1_adr1 = main_sram1_bus_adr1[8:0];
assign main_sram1_bus_dat_r1 = main_sram1_dat_r1;
assign main_sram1_dat_w = main_sram1_bus_dat_w1;

// synthesis translate_off
reg dummy_d_64;
// synthesis translate_on
always @(*) begin
	main_sram2_we <= 4'd0;
	main_sram2_we[0] <= (((main_sram2_bus_cyc1 & main_sram2_bus_stb1) & main_sram2_bus_we1) & main_sram2_bus_sel1[0]);
	main_sram2_we[1] <= (((main_sram2_bus_cyc1 & main_sram2_bus_stb1) & main_sram2_bus_we1) & main_sram2_bus_sel1[1]);
	main_sram2_we[2] <= (((main_sram2_bus_cyc1 & main_sram2_bus_stb1) & main_sram2_bus_we1) & main_sram2_bus_sel1[2]);
	main_sram2_we[3] <= (((main_sram2_bus_cyc1 & main_sram2_bus_stb1) & main_sram2_bus_we1) & main_sram2_bus_sel1[3]);
// synthesis translate_off
	dummy_d_64 <= dummy_s;
// synthesis translate_on
end
assign main_sram2_adr1 = main_sram2_bus_adr1[8:0];
assign main_sram2_bus_dat_r1 = main_sram2_dat_r1;
assign main_sram2_dat_w = main_sram2_bus_dat_w1;

// synthesis translate_off
reg dummy_d_65;
// synthesis translate_on
always @(*) begin
	main_sram3_we <= 4'd0;
	main_sram3_we[0] <= (((main_sram3_bus_cyc1 & main_sram3_bus_stb1) & main_sram3_bus_we1) & main_sram3_bus_sel1[0]);
	main_sram3_we[1] <= (((main_sram3_bus_cyc1 & main_sram3_bus_stb1) & main_sram3_bus_we1) & main_sram3_bus_sel1[1]);
	main_sram3_we[2] <= (((main_sram3_bus_cyc1 & main_sram3_bus_stb1) & main_sram3_bus_we1) & main_sram3_bus_sel1[2]);
	main_sram3_we[3] <= (((main_sram3_bus_cyc1 & main_sram3_bus_stb1) & main_sram3_bus_we1) & main_sram3_bus_sel1[3]);
// synthesis translate_off
	dummy_d_65 <= dummy_s;
// synthesis translate_on
end
assign main_sram3_adr1 = main_sram3_bus_adr1[8:0];
assign main_sram3_bus_dat_r1 = main_sram3_dat_r1;
assign main_sram3_dat_w = main_sram3_bus_dat_w1;

// synthesis translate_off
reg dummy_d_66;
// synthesis translate_on
always @(*) begin
	main_slave_sel <= 8'd0;
	main_slave_sel[0] <= (main_bus_adr[11:9] == 1'd0);
	main_slave_sel[1] <= (main_bus_adr[11:9] == 1'd1);
	main_slave_sel[2] <= (main_bus_adr[11:9] == 2'd2);
	main_slave_sel[3] <= (main_bus_adr[11:9] == 2'd3);
	main_slave_sel[4] <= (main_bus_adr[11:9] == 3'd4);
	main_slave_sel[5] <= (main_bus_adr[11:9] == 3'd5);
	main_slave_sel[6] <= (main_bus_adr[11:9] == 3'd6);
	main_slave_sel[7] <= (main_bus_adr[11:9] == 3'd7);
// synthesis translate_off
	dummy_d_66 <= dummy_s;
// synthesis translate_on
end
assign main_sram0_bus_adr0 = main_bus_adr;
assign main_sram0_bus_dat_w0 = main_bus_dat_w;
assign main_sram0_bus_sel0 = main_bus_sel;
assign main_sram0_bus_stb0 = main_bus_stb;
assign main_sram0_bus_we0 = main_bus_we;
assign main_sram0_bus_cti0 = main_bus_cti;
assign main_sram0_bus_bte0 = main_bus_bte;
assign main_sram1_bus_adr0 = main_bus_adr;
assign main_sram1_bus_dat_w0 = main_bus_dat_w;
assign main_sram1_bus_sel0 = main_bus_sel;
assign main_sram1_bus_stb0 = main_bus_stb;
assign main_sram1_bus_we0 = main_bus_we;
assign main_sram1_bus_cti0 = main_bus_cti;
assign main_sram1_bus_bte0 = main_bus_bte;
assign main_sram2_bus_adr0 = main_bus_adr;
assign main_sram2_bus_dat_w0 = main_bus_dat_w;
assign main_sram2_bus_sel0 = main_bus_sel;
assign main_sram2_bus_stb0 = main_bus_stb;
assign main_sram2_bus_we0 = main_bus_we;
assign main_sram2_bus_cti0 = main_bus_cti;
assign main_sram2_bus_bte0 = main_bus_bte;
assign main_sram3_bus_adr0 = main_bus_adr;
assign main_sram3_bus_dat_w0 = main_bus_dat_w;
assign main_sram3_bus_sel0 = main_bus_sel;
assign main_sram3_bus_stb0 = main_bus_stb;
assign main_sram3_bus_we0 = main_bus_we;
assign main_sram3_bus_cti0 = main_bus_cti;
assign main_sram3_bus_bte0 = main_bus_bte;
assign main_sram0_bus_adr1 = main_bus_adr;
assign main_sram0_bus_dat_w1 = main_bus_dat_w;
assign main_sram0_bus_sel1 = main_bus_sel;
assign main_sram0_bus_stb1 = main_bus_stb;
assign main_sram0_bus_we1 = main_bus_we;
assign main_sram0_bus_cti1 = main_bus_cti;
assign main_sram0_bus_bte1 = main_bus_bte;
assign main_sram1_bus_adr1 = main_bus_adr;
assign main_sram1_bus_dat_w1 = main_bus_dat_w;
assign main_sram1_bus_sel1 = main_bus_sel;
assign main_sram1_bus_stb1 = main_bus_stb;
assign main_sram1_bus_we1 = main_bus_we;
assign main_sram1_bus_cti1 = main_bus_cti;
assign main_sram1_bus_bte1 = main_bus_bte;
assign main_sram2_bus_adr1 = main_bus_adr;
assign main_sram2_bus_dat_w1 = main_bus_dat_w;
assign main_sram2_bus_sel1 = main_bus_sel;
assign main_sram2_bus_stb1 = main_bus_stb;
assign main_sram2_bus_we1 = main_bus_we;
assign main_sram2_bus_cti1 = main_bus_cti;
assign main_sram2_bus_bte1 = main_bus_bte;
assign main_sram3_bus_adr1 = main_bus_adr;
assign main_sram3_bus_dat_w1 = main_bus_dat_w;
assign main_sram3_bus_sel1 = main_bus_sel;
assign main_sram3_bus_stb1 = main_bus_stb;
assign main_sram3_bus_we1 = main_bus_we;
assign main_sram3_bus_cti1 = main_bus_cti;
assign main_sram3_bus_bte1 = main_bus_bte;
assign main_sram0_bus_cyc0 = (main_bus_cyc & main_slave_sel[0]);
assign main_sram1_bus_cyc0 = (main_bus_cyc & main_slave_sel[1]);
assign main_sram2_bus_cyc0 = (main_bus_cyc & main_slave_sel[2]);
assign main_sram3_bus_cyc0 = (main_bus_cyc & main_slave_sel[3]);
assign main_sram0_bus_cyc1 = (main_bus_cyc & main_slave_sel[4]);
assign main_sram1_bus_cyc1 = (main_bus_cyc & main_slave_sel[5]);
assign main_sram2_bus_cyc1 = (main_bus_cyc & main_slave_sel[6]);
assign main_sram3_bus_cyc1 = (main_bus_cyc & main_slave_sel[7]);
assign main_bus_ack = (((((((main_sram0_bus_ack0 | main_sram1_bus_ack0) | main_sram2_bus_ack0) | main_sram3_bus_ack0) | main_sram0_bus_ack1) | main_sram1_bus_ack1) | main_sram2_bus_ack1) | main_sram3_bus_ack1);
assign main_bus_err = (((((((main_sram0_bus_err0 | main_sram1_bus_err0) | main_sram2_bus_err0) | main_sram3_bus_err0) | main_sram0_bus_err1) | main_sram1_bus_err1) | main_sram2_bus_err1) | main_sram3_bus_err1);
assign main_bus_dat_r = (((((((({32{main_slave_sel_r[0]}} & main_sram0_bus_dat_r0) | ({32{main_slave_sel_r[1]}} & main_sram1_bus_dat_r0)) | ({32{main_slave_sel_r[2]}} & main_sram2_bus_dat_r0)) | ({32{main_slave_sel_r[3]}} & main_sram3_bus_dat_r0)) | ({32{main_slave_sel_r[4]}} & main_sram0_bus_dat_r1)) | ({32{main_slave_sel_r[5]}} & main_sram1_bus_dat_r1)) | ({32{main_slave_sel_r[6]}} & main_sram2_bus_dat_r1)) | ({32{main_slave_sel_r[7]}} & main_sram3_bus_dat_r1));
assign sys_kernel_clk = sys_clk;
assign sys_kernel_rst = main_kernel_cpu_storage;
assign main_kernel_cpu_ibus_adr = main_kernel_cpu_i_adr_o[31:2];
assign main_kernel_cpu_dbus_adr = main_kernel_cpu_d_adr_o[31:2];
assign builder_shared_adr = builder_comb_rhs_array_muxed0;
assign builder_shared_dat_w = builder_comb_rhs_array_muxed1;
assign builder_shared_sel = builder_comb_rhs_array_muxed2;
assign builder_shared_cyc = builder_comb_rhs_array_muxed3;
assign builder_shared_stb = builder_comb_rhs_array_muxed4;
assign builder_shared_we = builder_comb_rhs_array_muxed5;
assign builder_shared_cti = builder_comb_rhs_array_muxed6;
assign builder_shared_bte = builder_comb_rhs_array_muxed7;
assign main_kernel_cpu_ibus_dat_r = builder_shared_dat_r;
assign main_kernel_cpu_dbus_dat_r = builder_shared_dat_r;
assign main_kernel_cpu_ibus_ack = (builder_shared_ack & (builder_grant == 1'd0));
assign main_kernel_cpu_dbus_ack = (builder_shared_ack & (builder_grant == 1'd1));
assign main_kernel_cpu_ibus_err = (builder_shared_err & (builder_grant == 1'd0));
assign main_kernel_cpu_dbus_err = (builder_shared_err & (builder_grant == 1'd1));
assign builder_request = {(main_kernel_cpu_dbus_cyc & (~main_kernel_cpu_dbus_ack)), (main_kernel_cpu_ibus_cyc & (~main_kernel_cpu_ibus_ack))};

// synthesis translate_off
reg dummy_d_67;
// synthesis translate_on
always @(*) begin
	builder_slave_sel <= 5'd0;
	builder_slave_sel[0] <= ((1'd1 & (~builder_shared_adr[27])) & builder_shared_adr[28]);
	builder_slave_sel[1] <= ((1'd1 & builder_shared_adr[27]) & builder_shared_adr[28]);
	builder_slave_sel[2] <= (((1'd1 & (~builder_shared_adr[26])) & (~builder_shared_adr[28])) & builder_shared_adr[27]);
	builder_slave_sel[3] <= (((1'd1 & (~builder_shared_adr[28])) & builder_shared_adr[26]) & builder_shared_adr[27]);
	builder_slave_sel[4] <= ((1'd1 & (~builder_shared_adr[27])) & (~builder_shared_adr[28]));
// synthesis translate_off
	dummy_d_67 <= dummy_s;
// synthesis translate_on
end
assign main_kernel_cpu_wb_sdram_adr = builder_shared_adr;
assign main_kernel_cpu_wb_sdram_dat_w = builder_shared_dat_w;
assign main_kernel_cpu_wb_sdram_sel = builder_shared_sel;
assign main_kernel_cpu_wb_sdram_stb = builder_shared_stb;
assign main_kernel_cpu_wb_sdram_we = builder_shared_we;
assign main_kernel_cpu_wb_sdram_cti = builder_shared_cti;
assign main_kernel_cpu_wb_sdram_bte = builder_shared_bte;
assign main_mailbox_i2_adr = builder_shared_adr;
assign main_mailbox_i2_dat_w = builder_shared_dat_w;
assign main_mailbox_i2_sel = builder_shared_sel;
assign main_mailbox_i2_stb = builder_shared_stb;
assign main_mailbox_i2_we = builder_shared_we;
assign main_mailbox_i2_cti = builder_shared_cti;
assign main_mailbox_i2_bte = builder_shared_bte;
assign main_csrbank0_bus_adr = builder_shared_adr;
assign main_csrbank0_bus_dat_w = builder_shared_dat_w;
assign main_csrbank0_bus_sel = builder_shared_sel;
assign main_csrbank0_bus_stb = builder_shared_stb;
assign main_csrbank0_bus_we = builder_shared_we;
assign main_csrbank0_bus_cti = builder_shared_cti;
assign main_csrbank0_bus_bte = builder_shared_bte;
assign main_csrbank1_bus_adr = builder_shared_adr;
assign main_csrbank1_bus_dat_w = builder_shared_dat_w;
assign main_csrbank1_bus_sel = builder_shared_sel;
assign main_csrbank1_bus_stb = builder_shared_stb;
assign main_csrbank1_bus_we = builder_shared_we;
assign main_csrbank1_bus_cti = builder_shared_cti;
assign main_csrbank1_bus_bte = builder_shared_bte;
assign main_csrbank2_bus_adr = builder_shared_adr;
assign main_csrbank2_bus_dat_w = builder_shared_dat_w;
assign main_csrbank2_bus_sel = builder_shared_sel;
assign main_csrbank2_bus_stb = builder_shared_stb;
assign main_csrbank2_bus_we = builder_shared_we;
assign main_csrbank2_bus_cti = builder_shared_cti;
assign main_csrbank2_bus_bte = builder_shared_bte;
assign main_kernel_cpu_wb_sdram_cyc = (builder_shared_cyc & builder_slave_sel[0]);
assign main_mailbox_i2_cyc = (builder_shared_cyc & builder_slave_sel[1]);
assign main_csrbank0_bus_cyc = (builder_shared_cyc & builder_slave_sel[2]);
assign main_csrbank1_bus_cyc = (builder_shared_cyc & builder_slave_sel[3]);
assign main_csrbank2_bus_cyc = (builder_shared_cyc & builder_slave_sel[4]);
assign builder_shared_ack = ((((main_kernel_cpu_wb_sdram_ack | main_mailbox_i2_ack) | main_csrbank0_bus_ack) | main_csrbank1_bus_ack) | main_csrbank2_bus_ack);
assign builder_shared_err = ((((main_kernel_cpu_wb_sdram_err | main_mailbox_i2_err) | main_csrbank0_bus_err) | main_csrbank1_bus_err) | main_csrbank2_bus_err);
assign builder_shared_dat_r = ((((({32{builder_slave_sel_r[0]}} & main_kernel_cpu_wb_sdram_dat_r) | ({32{builder_slave_sel_r[1]}} & main_mailbox_i2_dat_r)) | ({32{builder_slave_sel_r[2]}} & main_csrbank0_bus_dat_r)) | ({32{builder_slave_sel_r[3]}} & main_csrbank1_bus_dat_r)) | ({32{builder_slave_sel_r[4]}} & main_csrbank2_bus_dat_r));
assign main_add_identifier_adr = main_add_identifier_storage;
assign main_add_identifier_status = main_add_identifier_dat_r;
assign main_zero_trigger = (main_value != 1'd0);
assign main_eventmanager_status_w = main_zero_status;

// synthesis translate_off
reg dummy_d_68;
// synthesis translate_on
always @(*) begin
	main_zero_clear <= 1'd0;
	if ((main_eventmanager_pending_re & main_eventmanager_pending_r)) begin
		main_zero_clear <= 1'd1;
	end
// synthesis translate_off
	dummy_d_68 <= dummy_s;
// synthesis translate_on
end
assign main_eventmanager_pending_w = main_zero_pending;
assign main_irq = (main_eventmanager_pending_w & main_eventmanager_storage);
assign main_zero_status = main_zero_trigger;
assign {user_led_1, user_led} = main_leds_storage;
assign main_i2c_tstriple0_o = main_i2c_out_storage[0];
assign main_i2c_tstriple0_oe = main_i2c_oe_storage[0];

// synthesis translate_off
reg dummy_d_69;
// synthesis translate_on
always @(*) begin
	main_i2c_status0 <= 2'd0;
	main_i2c_status0[0] <= main_i2c_status1;
	main_i2c_status0[1] <= main_i2c_status2;
// synthesis translate_off
	dummy_d_69 <= dummy_s;
// synthesis translate_on
end
assign main_i2c_tstriple1_o = main_i2c_out_storage[1];
assign main_i2c_tstriple1_oe = main_i2c_oe_storage[1];
assign ttl = main_output_8x0_pad_o;
assign ttl_1 = main_output_8x1_pad_o;
assign ttl_2 = main_output_8x2_pad_o;
assign main_inout_8x0_serdes_oe = main_inout_8x0_inout_8x0_oe;
assign main_inout_8x0_inout_8x0_input_state = main_inout_8x0_serdes_i0[7];
assign main_inout_8x0_inout_8x0_i = (main_inout_8x0_serdes_i0 ^ {8{main_inout_8x0_inout_8x0_i_d}});
assign main_inout_8x0_serdes_i0 = main_inout_8x0_serdes_i1;
assign main_inout_8x0_serdes_t_in = (~main_inout_8x0_serdes_oe);
assign main_inout_8x0_serdes_o1 = main_inout_8x0_serdes_o0;
assign main_inout_8x0_serdes_pad_i1 = main_inout_8x0_serdes_pad_i0;
assign main_inout_8x0_serdes_pad_o0 = main_inout_8x0_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_70;
// synthesis translate_on
always @(*) begin
	main_inout_8x0_inout_8x0_o <= 3'd0;
	if (main_inout_8x0_inout_8x0_i[7]) begin
		main_inout_8x0_inout_8x0_o <= 3'd7;
	end
	if (main_inout_8x0_inout_8x0_i[6]) begin
		main_inout_8x0_inout_8x0_o <= 3'd6;
	end
	if (main_inout_8x0_inout_8x0_i[5]) begin
		main_inout_8x0_inout_8x0_o <= 3'd5;
	end
	if (main_inout_8x0_inout_8x0_i[4]) begin
		main_inout_8x0_inout_8x0_o <= 3'd4;
	end
	if (main_inout_8x0_inout_8x0_i[3]) begin
		main_inout_8x0_inout_8x0_o <= 2'd3;
	end
	if (main_inout_8x0_inout_8x0_i[2]) begin
		main_inout_8x0_inout_8x0_o <= 2'd2;
	end
	if (main_inout_8x0_inout_8x0_i[1]) begin
		main_inout_8x0_inout_8x0_o <= 1'd1;
	end
	if (main_inout_8x0_inout_8x0_i[0]) begin
		main_inout_8x0_inout_8x0_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_70 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x0_inout_8x0_n = (main_inout_8x0_inout_8x0_i == 1'd0);
assign ttl_4 = main_output_8x3_pad_o;
assign ttl_5 = main_output_8x4_pad_o;
assign ttl_6 = main_output_8x5_pad_o;
assign main_inout_8x1_serdes_oe = main_inout_8x1_inout_8x1_oe;
assign main_inout_8x1_inout_8x1_input_state = main_inout_8x1_serdes_i0[7];
assign main_inout_8x1_inout_8x1_i = (main_inout_8x1_serdes_i0 ^ {8{main_inout_8x1_inout_8x1_i_d}});
assign main_inout_8x1_serdes_i0 = main_inout_8x1_serdes_i1;
assign main_inout_8x1_serdes_t_in = (~main_inout_8x1_serdes_oe);
assign main_inout_8x1_serdes_o1 = main_inout_8x1_serdes_o0;
assign main_inout_8x1_serdes_pad_i1 = main_inout_8x1_serdes_pad_i0;
assign main_inout_8x1_serdes_pad_o0 = main_inout_8x1_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_71;
// synthesis translate_on
always @(*) begin
	main_inout_8x1_inout_8x1_o <= 3'd0;
	if (main_inout_8x1_inout_8x1_i[7]) begin
		main_inout_8x1_inout_8x1_o <= 3'd7;
	end
	if (main_inout_8x1_inout_8x1_i[6]) begin
		main_inout_8x1_inout_8x1_o <= 3'd6;
	end
	if (main_inout_8x1_inout_8x1_i[5]) begin
		main_inout_8x1_inout_8x1_o <= 3'd5;
	end
	if (main_inout_8x1_inout_8x1_i[4]) begin
		main_inout_8x1_inout_8x1_o <= 3'd4;
	end
	if (main_inout_8x1_inout_8x1_i[3]) begin
		main_inout_8x1_inout_8x1_o <= 2'd3;
	end
	if (main_inout_8x1_inout_8x1_i[2]) begin
		main_inout_8x1_inout_8x1_o <= 2'd2;
	end
	if (main_inout_8x1_inout_8x1_i[1]) begin
		main_inout_8x1_inout_8x1_o <= 1'd1;
	end
	if (main_inout_8x1_inout_8x1_i[0]) begin
		main_inout_8x1_inout_8x1_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_71 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x1_inout_8x1_n = (main_inout_8x1_inout_8x1_i == 1'd0);
assign ttl_8 = main_output_8x6_pad_o;
assign ttl_9 = main_output_8x7_pad_o;
assign ttl_10 = main_output_8x8_pad_o;
assign main_inout_8x2_serdes_oe = main_inout_8x2_inout_8x2_oe;
assign main_inout_8x2_inout_8x2_input_state = main_inout_8x2_serdes_i0[7];
assign main_inout_8x2_inout_8x2_i = (main_inout_8x2_serdes_i0 ^ {8{main_inout_8x2_inout_8x2_i_d}});
assign main_inout_8x2_serdes_i0 = main_inout_8x2_serdes_i1;
assign main_inout_8x2_serdes_t_in = (~main_inout_8x2_serdes_oe);
assign main_inout_8x2_serdes_o1 = main_inout_8x2_serdes_o0;
assign main_inout_8x2_serdes_pad_i1 = main_inout_8x2_serdes_pad_i0;
assign main_inout_8x2_serdes_pad_o0 = main_inout_8x2_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_72;
// synthesis translate_on
always @(*) begin
	main_inout_8x2_inout_8x2_o <= 3'd0;
	if (main_inout_8x2_inout_8x2_i[7]) begin
		main_inout_8x2_inout_8x2_o <= 3'd7;
	end
	if (main_inout_8x2_inout_8x2_i[6]) begin
		main_inout_8x2_inout_8x2_o <= 3'd6;
	end
	if (main_inout_8x2_inout_8x2_i[5]) begin
		main_inout_8x2_inout_8x2_o <= 3'd5;
	end
	if (main_inout_8x2_inout_8x2_i[4]) begin
		main_inout_8x2_inout_8x2_o <= 3'd4;
	end
	if (main_inout_8x2_inout_8x2_i[3]) begin
		main_inout_8x2_inout_8x2_o <= 2'd3;
	end
	if (main_inout_8x2_inout_8x2_i[2]) begin
		main_inout_8x2_inout_8x2_o <= 2'd2;
	end
	if (main_inout_8x2_inout_8x2_i[1]) begin
		main_inout_8x2_inout_8x2_o <= 1'd1;
	end
	if (main_inout_8x2_inout_8x2_i[0]) begin
		main_inout_8x2_inout_8x2_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_72 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x2_inout_8x2_n = (main_inout_8x2_inout_8x2_i == 1'd0);
assign ttl_12 = main_output_8x9_pad_o;
assign ttl_13 = main_output_8x10_pad_o;
assign ttl_14 = main_output_8x11_pad_o;
assign main_inout_8x3_serdes_oe = main_inout_8x3_inout_8x3_oe;
assign main_inout_8x3_inout_8x3_input_state = main_inout_8x3_serdes_i0[7];
assign main_inout_8x3_inout_8x3_i = (main_inout_8x3_serdes_i0 ^ {8{main_inout_8x3_inout_8x3_i_d}});
assign main_inout_8x3_serdes_i0 = main_inout_8x3_serdes_i1;
assign main_inout_8x3_serdes_t_in = (~main_inout_8x3_serdes_oe);
assign main_inout_8x3_serdes_o1 = main_inout_8x3_serdes_o0;
assign main_inout_8x3_serdes_pad_i1 = main_inout_8x3_serdes_pad_i0;
assign main_inout_8x3_serdes_pad_o0 = main_inout_8x3_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_73;
// synthesis translate_on
always @(*) begin
	main_inout_8x3_inout_8x3_o <= 3'd0;
	if (main_inout_8x3_inout_8x3_i[7]) begin
		main_inout_8x3_inout_8x3_o <= 3'd7;
	end
	if (main_inout_8x3_inout_8x3_i[6]) begin
		main_inout_8x3_inout_8x3_o <= 3'd6;
	end
	if (main_inout_8x3_inout_8x3_i[5]) begin
		main_inout_8x3_inout_8x3_o <= 3'd5;
	end
	if (main_inout_8x3_inout_8x3_i[4]) begin
		main_inout_8x3_inout_8x3_o <= 3'd4;
	end
	if (main_inout_8x3_inout_8x3_i[3]) begin
		main_inout_8x3_inout_8x3_o <= 2'd3;
	end
	if (main_inout_8x3_inout_8x3_i[2]) begin
		main_inout_8x3_inout_8x3_o <= 2'd2;
	end
	if (main_inout_8x3_inout_8x3_i[1]) begin
		main_inout_8x3_inout_8x3_o <= 1'd1;
	end
	if (main_inout_8x3_inout_8x3_i[0]) begin
		main_inout_8x3_inout_8x3_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_73 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x3_inout_8x3_n = (main_inout_8x3_inout_8x3_i == 1'd0);
assign main_inout_8x4_serdes_oe = main_inout_8x4_inout_8x4_oe;
assign main_inout_8x4_inout_8x4_input_state = main_inout_8x4_serdes_i0[7];
assign main_inout_8x4_inout_8x4_i = (main_inout_8x4_serdes_i0 ^ {8{main_inout_8x4_inout_8x4_i_d}});
assign main_inout_8x4_serdes_i0 = main_inout_8x4_serdes_i1;
assign main_inout_8x4_serdes_t_in = (~main_inout_8x4_serdes_oe);
assign main_inout_8x4_serdes_o1 = main_inout_8x4_serdes_o0;
assign main_inout_8x4_serdes_pad_i1 = main_inout_8x4_serdes_pad_i0;
assign main_inout_8x4_serdes_pad_o0 = main_inout_8x4_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_74;
// synthesis translate_on
always @(*) begin
	main_inout_8x4_inout_8x4_o <= 3'd0;
	if (main_inout_8x4_inout_8x4_i[7]) begin
		main_inout_8x4_inout_8x4_o <= 3'd7;
	end
	if (main_inout_8x4_inout_8x4_i[6]) begin
		main_inout_8x4_inout_8x4_o <= 3'd6;
	end
	if (main_inout_8x4_inout_8x4_i[5]) begin
		main_inout_8x4_inout_8x4_o <= 3'd5;
	end
	if (main_inout_8x4_inout_8x4_i[4]) begin
		main_inout_8x4_inout_8x4_o <= 3'd4;
	end
	if (main_inout_8x4_inout_8x4_i[3]) begin
		main_inout_8x4_inout_8x4_o <= 2'd3;
	end
	if (main_inout_8x4_inout_8x4_i[2]) begin
		main_inout_8x4_inout_8x4_o <= 2'd2;
	end
	if (main_inout_8x4_inout_8x4_i[1]) begin
		main_inout_8x4_inout_8x4_o <= 1'd1;
	end
	if (main_inout_8x4_inout_8x4_i[0]) begin
		main_inout_8x4_inout_8x4_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_74 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x4_inout_8x4_n = (main_inout_8x4_inout_8x4_i == 1'd0);
assign main_inout_8x5_serdes_oe = main_inout_8x5_inout_8x5_oe;
assign main_inout_8x5_inout_8x5_input_state = main_inout_8x5_serdes_i0[7];
assign main_inout_8x5_inout_8x5_i = (main_inout_8x5_serdes_i0 ^ {8{main_inout_8x5_inout_8x5_i_d}});
assign main_inout_8x5_serdes_i0 = main_inout_8x5_serdes_i1;
assign main_inout_8x5_serdes_t_in = (~main_inout_8x5_serdes_oe);
assign main_inout_8x5_serdes_o1 = main_inout_8x5_serdes_o0;
assign main_inout_8x5_serdes_pad_i1 = main_inout_8x5_serdes_pad_i0;
assign main_inout_8x5_serdes_pad_o0 = main_inout_8x5_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_75;
// synthesis translate_on
always @(*) begin
	main_inout_8x5_inout_8x5_o <= 3'd0;
	if (main_inout_8x5_inout_8x5_i[7]) begin
		main_inout_8x5_inout_8x5_o <= 3'd7;
	end
	if (main_inout_8x5_inout_8x5_i[6]) begin
		main_inout_8x5_inout_8x5_o <= 3'd6;
	end
	if (main_inout_8x5_inout_8x5_i[5]) begin
		main_inout_8x5_inout_8x5_o <= 3'd5;
	end
	if (main_inout_8x5_inout_8x5_i[4]) begin
		main_inout_8x5_inout_8x5_o <= 3'd4;
	end
	if (main_inout_8x5_inout_8x5_i[3]) begin
		main_inout_8x5_inout_8x5_o <= 2'd3;
	end
	if (main_inout_8x5_inout_8x5_i[2]) begin
		main_inout_8x5_inout_8x5_o <= 2'd2;
	end
	if (main_inout_8x5_inout_8x5_i[1]) begin
		main_inout_8x5_inout_8x5_o <= 1'd1;
	end
	if (main_inout_8x5_inout_8x5_i[0]) begin
		main_inout_8x5_inout_8x5_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_75 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x5_inout_8x5_n = (main_inout_8x5_inout_8x5_i == 1'd0);
assign main_inout_8x6_serdes_oe = main_inout_8x6_inout_8x6_oe;
assign main_inout_8x6_inout_8x6_input_state = main_inout_8x6_serdes_i0[7];
assign main_inout_8x6_inout_8x6_i = (main_inout_8x6_serdes_i0 ^ {8{main_inout_8x6_inout_8x6_i_d}});
assign main_inout_8x6_serdes_i0 = main_inout_8x6_serdes_i1;
assign main_inout_8x6_serdes_t_in = (~main_inout_8x6_serdes_oe);
assign main_inout_8x6_serdes_o1 = main_inout_8x6_serdes_o0;
assign main_inout_8x6_serdes_pad_i1 = main_inout_8x6_serdes_pad_i0;
assign main_inout_8x6_serdes_pad_o0 = main_inout_8x6_serdes_pad_o1;

// synthesis translate_off
reg dummy_d_76;
// synthesis translate_on
always @(*) begin
	main_inout_8x6_inout_8x6_o <= 3'd0;
	if (main_inout_8x6_inout_8x6_i[7]) begin
		main_inout_8x6_inout_8x6_o <= 3'd7;
	end
	if (main_inout_8x6_inout_8x6_i[6]) begin
		main_inout_8x6_inout_8x6_o <= 3'd6;
	end
	if (main_inout_8x6_inout_8x6_i[5]) begin
		main_inout_8x6_inout_8x6_o <= 3'd5;
	end
	if (main_inout_8x6_inout_8x6_i[4]) begin
		main_inout_8x6_inout_8x6_o <= 3'd4;
	end
	if (main_inout_8x6_inout_8x6_i[3]) begin
		main_inout_8x6_inout_8x6_o <= 2'd3;
	end
	if (main_inout_8x6_inout_8x6_i[2]) begin
		main_inout_8x6_inout_8x6_o <= 2'd2;
	end
	if (main_inout_8x6_inout_8x6_i[1]) begin
		main_inout_8x6_inout_8x6_o <= 1'd1;
	end
	if (main_inout_8x6_inout_8x6_i[0]) begin
		main_inout_8x6_inout_8x6_o <= 1'd0;
	end
// synthesis translate_off
	dummy_d_76 <= dummy_s;
// synthesis translate_on
end
assign main_inout_8x6_inout_8x6_n = (main_inout_8x6_inout_8x6_i == 1'd0);
assign user_led_2 = main_output0_pad_o;
assign ams101_dac_ldac = main_output1_pad_o;
assign main_spimaster0_spimachine0_length = main_spimaster0_config_length;
assign main_spimaster0_spimachine0_end0 = main_spimaster0_config_end;
assign main_spimaster0_spimachine0_div = main_spimaster0_config_div;
assign main_spimaster0_spimachine0_clk_phase = main_spimaster0_config_clk_phase;
assign main_spimaster0_spimachine0_lsb_first = main_spimaster0_config_lsb_first;
assign main_spimaster0_interface_half_duplex = main_spimaster0_config_half_duplex;
assign main_spimaster0_interface_cs = main_spimaster0_config_cs;
assign main_spimaster0_interface_cs_polarity = {1{main_spimaster0_config_cs_polarity}};
assign main_spimaster0_interface_clk_polarity = main_spimaster0_config_clk_polarity;
assign main_spimaster0_interface_offline = main_spimaster0_config_offline;
assign main_spimaster0_interface_cs_next = main_spimaster0_spimachine0_cs_next;
assign main_spimaster0_interface_clk_next = main_spimaster0_spimachine0_clk_next;
assign main_spimaster0_interface_ce = main_spimaster0_spimachine0_ce;
assign main_spimaster0_interface_sample = main_spimaster0_spimachine0_sample;
assign main_spimaster0_spimachine0_sdi = main_spimaster0_interface_sdi;
assign main_spimaster0_interface_sdo = main_spimaster0_spimachine0_sdo;
assign main_spimaster0_spimachine0_load0 = ((main_spimaster0_ointerface0_stb & main_spimaster0_spimachine0_writable) & (~main_spimaster0_ointerface0_address));
assign main_spimaster0_spimachine0_pdo = main_spimaster0_ointerface0_data;
assign main_spimaster0_ointerface0_busy = (~main_spimaster0_spimachine0_writable);
assign main_spimaster0_iinterface0_stb = (main_spimaster0_spimachine0_readable & main_spimaster0_read);
assign main_spimaster0_iinterface0_data = main_spimaster0_spimachine0_pdi;
assign main_spimaster0_interface_miso_oe = 1'd0;
assign main_spimaster0_interface_mosi_o = main_spimaster0_interface_sdo;
assign main_spimaster0_interface_miso_o = main_spimaster0_interface_sdo;
assign main_spimaster0_interface_cs_oe = (~main_spimaster0_interface_offline);
assign main_spimaster0_interface_clk_oe = (~main_spimaster0_interface_offline);
assign main_spimaster0_interface_mosi_oe = (~(main_spimaster0_interface_offline | main_spimaster0_interface_half_duplex));

// synthesis translate_off
reg dummy_d_77;
// synthesis translate_on
always @(*) begin
	main_spimaster0_interface_sdi <= 1'd0;
	if ((main_spimaster0_interface_cs != 1'd0)) begin
		main_spimaster0_interface_sdi <= (main_spimaster0_interface_half_duplex ? main_spimaster0_interface_mosi_reg : main_spimaster0_interface_miso_reg);
	end
// synthesis translate_off
	dummy_d_77 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster0_spimachine0_ce = (main_spimaster0_spimachine0_done & main_spimaster0_spimachine0_count);
assign main_spimaster0_spimachine0_pdi = (main_spimaster0_spimachine0_lsb_first ? {main_spimaster0_spimachine0_sdi, main_spimaster0_spimachine0_sr[31:1]} : {main_spimaster0_spimachine0_sr[30:0], main_spimaster0_spimachine0_sdi});
assign main_spimaster0_spimachine0_cnt_done = (main_spimaster0_spimachine0_cnt == 1'd0);
assign main_spimaster0_spimachine0_done = (main_spimaster0_spimachine0_cnt_done & (~main_spimaster0_spimachine0_do_extend));

// synthesis translate_off
reg dummy_d_78;
// synthesis translate_on
always @(*) begin
	main_spimaster0_spimachine0_clk_next <= 1'd0;
	main_spimaster0_spimachine0_cs_next <= 1'd0;
	main_spimaster0_spimachine0_idle <= 1'd0;
	main_spimaster0_spimachine0_readable <= 1'd0;
	main_spimaster0_spimachine0_writable <= 1'd0;
	main_spimaster0_spimachine0_load1 <= 1'd0;
	main_spimaster0_spimachine0_shift <= 1'd0;
	main_spimaster0_spimachine0_sample <= 1'd0;
	main_spimaster0_spimachine0_extend <= 1'd0;
	main_spimaster0_spimachine0_count <= 1'd0;
	builder_spimaster0_next_state <= 3'd0;
	builder_spimaster0_next_state <= builder_spimaster0_state;
	case (builder_spimaster0_state)
		1'd1: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_extend <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= 1'd1;
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= (~main_spimaster0_spimachine0_clk_phase);
			if (main_spimaster0_spimachine0_done) begin
				main_spimaster0_spimachine0_sample <= 1'd1;
				builder_spimaster0_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			main_spimaster0_spimachine0_count <= 1'd1;
			main_spimaster0_spimachine0_extend <= 1'd1;
			main_spimaster0_spimachine0_clk_next <= main_spimaster0_spimachine0_clk_phase;
			if (main_spimaster0_spimachine0_done) begin
				if ((main_spimaster0_spimachine0_n == 1'd0)) begin
					main_spimaster0_spimachine0_readable <= 1'd1;
					main_spimaster0_spimachine0_writable <= 1'd1;
					if (main_spimaster0_spimachine0_end1) begin
						main_spimaster0_spimachine0_clk_next <= 1'd0;
						main_spimaster0_spimachine0_writable <= 1'd0;
						if (main_spimaster0_spimachine0_clk_phase) begin
							main_spimaster0_spimachine0_cs_next <= 1'd0;
							builder_spimaster0_next_state <= 3'd5;
						end else begin
							builder_spimaster0_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster0_spimachine0_load0) begin
							main_spimaster0_spimachine0_load1 <= 1'd1;
							builder_spimaster0_next_state <= 2'd2;
						end else begin
							main_spimaster0_spimachine0_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster0_spimachine0_shift <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster0_spimachine0_count <= 1'd1;
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster0_spimachine0_done) begin
				builder_spimaster0_next_state <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster0_spimachine0_idle <= 1'd1;
			main_spimaster0_spimachine0_writable <= 1'd1;
			main_spimaster0_spimachine0_cs_next <= 1'd1;
			if (main_spimaster0_spimachine0_load0) begin
				main_spimaster0_spimachine0_count <= 1'd1;
				main_spimaster0_spimachine0_load1 <= 1'd1;
				if (main_spimaster0_spimachine0_clk_phase) begin
					builder_spimaster0_next_state <= 1'd1;
				end else begin
					main_spimaster0_spimachine0_extend <= 1'd1;
					builder_spimaster0_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_78 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster1_spimachine1_length = main_spimaster1_config_length;
assign main_spimaster1_spimachine1_end0 = main_spimaster1_config_end;
assign main_spimaster1_spimachine1_div = main_spimaster1_config_div;
assign main_spimaster1_spimachine1_clk_phase = main_spimaster1_config_clk_phase;
assign main_spimaster1_spimachine1_lsb_first = main_spimaster1_config_lsb_first;
assign main_spimaster1_interface_half_duplex = main_spimaster1_config_half_duplex;
assign main_spimaster1_interface_cs = main_spimaster1_config_cs;
assign main_spimaster1_interface_cs_polarity = {1{main_spimaster1_config_cs_polarity}};
assign main_spimaster1_interface_clk_polarity = main_spimaster1_config_clk_polarity;
assign main_spimaster1_interface_offline = main_spimaster1_config_offline;
assign main_spimaster1_interface_cs_next = main_spimaster1_spimachine1_cs_next;
assign main_spimaster1_interface_clk_next = main_spimaster1_spimachine1_clk_next;
assign main_spimaster1_interface_ce = main_spimaster1_spimachine1_ce;
assign main_spimaster1_interface_sample = main_spimaster1_spimachine1_sample;
assign main_spimaster1_spimachine1_sdi = main_spimaster1_interface_sdi;
assign main_spimaster1_interface_sdo = main_spimaster1_spimachine1_sdo;
assign main_spimaster1_spimachine1_load0 = ((main_spimaster1_ointerface1_stb & main_spimaster1_spimachine1_writable) & (~main_spimaster1_ointerface1_address));
assign main_spimaster1_spimachine1_pdo = main_spimaster1_ointerface1_data;
assign main_spimaster1_ointerface1_busy = (~main_spimaster1_spimachine1_writable);
assign main_spimaster1_iinterface1_stb = (main_spimaster1_spimachine1_readable & main_spimaster1_read);
assign main_spimaster1_iinterface1_data = main_spimaster1_spimachine1_pdi;
assign main_spimaster1_interface_miso_oe = 1'd0;
assign main_spimaster1_interface_mosi_o = main_spimaster1_interface_sdo;
assign main_spimaster1_interface_miso_o = main_spimaster1_interface_sdo;
assign main_spimaster1_interface_cs_oe = (~main_spimaster1_interface_offline);
assign main_spimaster1_interface_clk_oe = (~main_spimaster1_interface_offline);
assign main_spimaster1_interface_mosi_oe = (~(main_spimaster1_interface_offline | main_spimaster1_interface_half_duplex));

// synthesis translate_off
reg dummy_d_79;
// synthesis translate_on
always @(*) begin
	main_spimaster1_interface_sdi <= 1'd0;
	if ((main_spimaster1_interface_cs != 1'd0)) begin
		main_spimaster1_interface_sdi <= (main_spimaster1_interface_half_duplex ? main_spimaster1_interface_mosi_reg : main_spimaster1_interface_miso_reg);
	end
// synthesis translate_off
	dummy_d_79 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster1_spimachine1_ce = (main_spimaster1_spimachine1_done & main_spimaster1_spimachine1_count);
assign main_spimaster1_spimachine1_pdi = (main_spimaster1_spimachine1_lsb_first ? {main_spimaster1_spimachine1_sdi, main_spimaster1_spimachine1_sr[31:1]} : {main_spimaster1_spimachine1_sr[30:0], main_spimaster1_spimachine1_sdi});
assign main_spimaster1_spimachine1_cnt_done = (main_spimaster1_spimachine1_cnt == 1'd0);
assign main_spimaster1_spimachine1_done = (main_spimaster1_spimachine1_cnt_done & (~main_spimaster1_spimachine1_do_extend));

// synthesis translate_off
reg dummy_d_80;
// synthesis translate_on
always @(*) begin
	main_spimaster1_spimachine1_clk_next <= 1'd0;
	main_spimaster1_spimachine1_cs_next <= 1'd0;
	main_spimaster1_spimachine1_idle <= 1'd0;
	main_spimaster1_spimachine1_readable <= 1'd0;
	main_spimaster1_spimachine1_writable <= 1'd0;
	main_spimaster1_spimachine1_load1 <= 1'd0;
	main_spimaster1_spimachine1_shift <= 1'd0;
	main_spimaster1_spimachine1_sample <= 1'd0;
	main_spimaster1_spimachine1_extend <= 1'd0;
	main_spimaster1_spimachine1_count <= 1'd0;
	builder_spimaster1_next_state <= 3'd0;
	builder_spimaster1_next_state <= builder_spimaster1_state;
	case (builder_spimaster1_state)
		1'd1: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_extend <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= 1'd1;
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= (~main_spimaster1_spimachine1_clk_phase);
			if (main_spimaster1_spimachine1_done) begin
				main_spimaster1_spimachine1_sample <= 1'd1;
				builder_spimaster1_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			main_spimaster1_spimachine1_count <= 1'd1;
			main_spimaster1_spimachine1_extend <= 1'd1;
			main_spimaster1_spimachine1_clk_next <= main_spimaster1_spimachine1_clk_phase;
			if (main_spimaster1_spimachine1_done) begin
				if ((main_spimaster1_spimachine1_n == 1'd0)) begin
					main_spimaster1_spimachine1_readable <= 1'd1;
					main_spimaster1_spimachine1_writable <= 1'd1;
					if (main_spimaster1_spimachine1_end1) begin
						main_spimaster1_spimachine1_clk_next <= 1'd0;
						main_spimaster1_spimachine1_writable <= 1'd0;
						if (main_spimaster1_spimachine1_clk_phase) begin
							main_spimaster1_spimachine1_cs_next <= 1'd0;
							builder_spimaster1_next_state <= 3'd5;
						end else begin
							builder_spimaster1_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster1_spimachine1_load0) begin
							main_spimaster1_spimachine1_load1 <= 1'd1;
							builder_spimaster1_next_state <= 2'd2;
						end else begin
							main_spimaster1_spimachine1_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster1_spimachine1_shift <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster1_spimachine1_count <= 1'd1;
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster1_spimachine1_done) begin
				builder_spimaster1_next_state <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster1_spimachine1_idle <= 1'd1;
			main_spimaster1_spimachine1_writable <= 1'd1;
			main_spimaster1_spimachine1_cs_next <= 1'd1;
			if (main_spimaster1_spimachine1_load0) begin
				main_spimaster1_spimachine1_count <= 1'd1;
				main_spimaster1_spimachine1_load1 <= 1'd1;
				if (main_spimaster1_spimachine1_clk_phase) begin
					builder_spimaster1_next_state <= 1'd1;
				end else begin
					main_spimaster1_spimachine1_extend <= 1'd1;
					builder_spimaster1_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_80 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster2_spimachine2_length = main_spimaster2_config_length;
assign main_spimaster2_spimachine2_end0 = main_spimaster2_config_end;
assign main_spimaster2_spimachine2_div = main_spimaster2_config_div;
assign main_spimaster2_spimachine2_clk_phase = main_spimaster2_config_clk_phase;
assign main_spimaster2_spimachine2_lsb_first = main_spimaster2_config_lsb_first;
assign main_spimaster2_interface_half_duplex = main_spimaster2_config_half_duplex;
assign main_spimaster2_interface_cs = main_spimaster2_config_cs;
assign main_spimaster2_interface_cs_polarity = {1{main_spimaster2_config_cs_polarity}};
assign main_spimaster2_interface_clk_polarity = main_spimaster2_config_clk_polarity;
assign main_spimaster2_interface_offline = main_spimaster2_config_offline;
assign main_spimaster2_interface_cs_next = main_spimaster2_spimachine2_cs_next;
assign main_spimaster2_interface_clk_next = main_spimaster2_spimachine2_clk_next;
assign main_spimaster2_interface_ce = main_spimaster2_spimachine2_ce;
assign main_spimaster2_interface_sample = main_spimaster2_spimachine2_sample;
assign main_spimaster2_spimachine2_sdi = main_spimaster2_interface_sdi;
assign main_spimaster2_interface_sdo = main_spimaster2_spimachine2_sdo;
assign main_spimaster2_spimachine2_load0 = ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable) & (~main_spimaster2_ointerface2_address));
assign main_spimaster2_spimachine2_pdo = main_spimaster2_ointerface2_data;
assign main_spimaster2_ointerface2_busy = (~main_spimaster2_spimachine2_writable);
assign main_spimaster2_iinterface2_stb = (main_spimaster2_spimachine2_readable & main_spimaster2_read);
assign main_spimaster2_iinterface2_data = main_spimaster2_spimachine2_pdi;
assign main_spimaster2_interface_miso_oe = 1'd0;
assign main_spimaster2_interface_mosi_o = main_spimaster2_interface_sdo;
assign main_spimaster2_interface_miso_o = main_spimaster2_interface_sdo;
assign main_spimaster2_interface_cs_oe = (~main_spimaster2_interface_offline);
assign main_spimaster2_interface_clk_oe = (~main_spimaster2_interface_offline);
assign main_spimaster2_interface_mosi_oe = (~(main_spimaster2_interface_offline | main_spimaster2_interface_half_duplex));

// synthesis translate_off
reg dummy_d_81;
// synthesis translate_on
always @(*) begin
	main_spimaster2_interface_sdi <= 1'd0;
	if ((main_spimaster2_interface_cs != 1'd0)) begin
		main_spimaster2_interface_sdi <= (main_spimaster2_interface_half_duplex ? main_spimaster2_interface_mosi_reg : main_spimaster2_interface_miso_reg);
	end
// synthesis translate_off
	dummy_d_81 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster2_spimachine2_ce = (main_spimaster2_spimachine2_done & main_spimaster2_spimachine2_count);
assign main_spimaster2_spimachine2_pdi = (main_spimaster2_spimachine2_lsb_first ? {main_spimaster2_spimachine2_sdi, main_spimaster2_spimachine2_sr[31:1]} : {main_spimaster2_spimachine2_sr[30:0], main_spimaster2_spimachine2_sdi});
assign main_spimaster2_spimachine2_cnt_done = (main_spimaster2_spimachine2_cnt == 1'd0);
assign main_spimaster2_spimachine2_done = (main_spimaster2_spimachine2_cnt_done & (~main_spimaster2_spimachine2_do_extend));

// synthesis translate_off
reg dummy_d_82;
// synthesis translate_on
always @(*) begin
	main_spimaster2_spimachine2_clk_next <= 1'd0;
	main_spimaster2_spimachine2_cs_next <= 1'd0;
	main_spimaster2_spimachine2_idle <= 1'd0;
	main_spimaster2_spimachine2_readable <= 1'd0;
	main_spimaster2_spimachine2_writable <= 1'd0;
	main_spimaster2_spimachine2_load1 <= 1'd0;
	main_spimaster2_spimachine2_shift <= 1'd0;
	main_spimaster2_spimachine2_sample <= 1'd0;
	main_spimaster2_spimachine2_extend <= 1'd0;
	main_spimaster2_spimachine2_count <= 1'd0;
	builder_spimaster2_next_state <= 3'd0;
	builder_spimaster2_next_state <= builder_spimaster2_state;
	case (builder_spimaster2_state)
		1'd1: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= (~main_spimaster2_spimachine2_clk_phase);
			if (main_spimaster2_spimachine2_done) begin
				main_spimaster2_spimachine2_sample <= 1'd1;
				builder_spimaster2_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			main_spimaster2_spimachine2_count <= 1'd1;
			main_spimaster2_spimachine2_extend <= 1'd1;
			main_spimaster2_spimachine2_clk_next <= main_spimaster2_spimachine2_clk_phase;
			if (main_spimaster2_spimachine2_done) begin
				if ((main_spimaster2_spimachine2_n == 1'd0)) begin
					main_spimaster2_spimachine2_readable <= 1'd1;
					main_spimaster2_spimachine2_writable <= 1'd1;
					if (main_spimaster2_spimachine2_end1) begin
						main_spimaster2_spimachine2_clk_next <= 1'd0;
						main_spimaster2_spimachine2_writable <= 1'd0;
						if (main_spimaster2_spimachine2_clk_phase) begin
							main_spimaster2_spimachine2_cs_next <= 1'd0;
							builder_spimaster2_next_state <= 3'd5;
						end else begin
							builder_spimaster2_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster2_spimachine2_load0) begin
							main_spimaster2_spimachine2_load1 <= 1'd1;
							builder_spimaster2_next_state <= 2'd2;
						end else begin
							main_spimaster2_spimachine2_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster2_spimachine2_shift <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster2_spimachine2_count <= 1'd1;
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster2_spimachine2_done) begin
				builder_spimaster2_next_state <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster2_spimachine2_idle <= 1'd1;
			main_spimaster2_spimachine2_writable <= 1'd1;
			main_spimaster2_spimachine2_cs_next <= 1'd1;
			if (main_spimaster2_spimachine2_load0) begin
				main_spimaster2_spimachine2_count <= 1'd1;
				main_spimaster2_spimachine2_load1 <= 1'd1;
				if (main_spimaster2_spimachine2_clk_phase) begin
					builder_spimaster2_next_state <= 1'd1;
				end else begin
					main_spimaster2_spimachine2_extend <= 1'd1;
					builder_spimaster2_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_82 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster3_spimachine3_length = main_spimaster3_config_length;
assign main_spimaster3_spimachine3_end0 = main_spimaster3_config_end;
assign main_spimaster3_spimachine3_div = main_spimaster3_config_div;
assign main_spimaster3_spimachine3_clk_phase = main_spimaster3_config_clk_phase;
assign main_spimaster3_spimachine3_lsb_first = main_spimaster3_config_lsb_first;
assign main_spimaster3_interface_half_duplex = main_spimaster3_config_half_duplex;
assign main_spimaster3_interface_cs = main_spimaster3_config_cs;
assign main_spimaster3_interface_cs_polarity = {1{main_spimaster3_config_cs_polarity}};
assign main_spimaster3_interface_clk_polarity = main_spimaster3_config_clk_polarity;
assign main_spimaster3_interface_offline = main_spimaster3_config_offline;
assign main_spimaster3_interface_cs_next = main_spimaster3_spimachine3_cs_next;
assign main_spimaster3_interface_clk_next = main_spimaster3_spimachine3_clk_next;
assign main_spimaster3_interface_ce = main_spimaster3_spimachine3_ce;
assign main_spimaster3_interface_sample = main_spimaster3_spimachine3_sample;
assign main_spimaster3_spimachine3_sdi = main_spimaster3_interface_sdi;
assign main_spimaster3_interface_sdo = main_spimaster3_spimachine3_sdo;
assign main_spimaster3_spimachine3_load0 = ((main_spimaster3_ointerface3_stb & main_spimaster3_spimachine3_writable) & (~main_spimaster3_ointerface3_address));
assign main_spimaster3_spimachine3_pdo = main_spimaster3_ointerface3_data;
assign main_spimaster3_ointerface3_busy = (~main_spimaster3_spimachine3_writable);
assign main_spimaster3_iinterface3_stb = (main_spimaster3_spimachine3_readable & main_spimaster3_read);
assign main_spimaster3_iinterface3_data = main_spimaster3_spimachine3_pdi;
assign main_spimaster3_interface_miso_oe = 1'd0;
assign main_spimaster3_interface_mosi_o = main_spimaster3_interface_sdo;
assign main_spimaster3_interface_miso_o = main_spimaster3_interface_sdo;
assign main_spimaster3_interface_cs_oe = (~main_spimaster3_interface_offline);
assign main_spimaster3_interface_clk_oe = (~main_spimaster3_interface_offline);
assign main_spimaster3_interface_mosi_oe = (~(main_spimaster3_interface_offline | main_spimaster3_interface_half_duplex));

// synthesis translate_off
reg dummy_d_83;
// synthesis translate_on
always @(*) begin
	main_spimaster3_interface_sdi <= 1'd0;
	if ((main_spimaster3_interface_cs != 1'd0)) begin
		main_spimaster3_interface_sdi <= (main_spimaster3_interface_half_duplex ? main_spimaster3_interface_mosi_reg : main_spimaster3_interface_miso_reg);
	end
// synthesis translate_off
	dummy_d_83 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster3_spimachine3_ce = (main_spimaster3_spimachine3_done & main_spimaster3_spimachine3_count);
assign main_spimaster3_spimachine3_pdi = (main_spimaster3_spimachine3_lsb_first ? {main_spimaster3_spimachine3_sdi, main_spimaster3_spimachine3_sr[31:1]} : {main_spimaster3_spimachine3_sr[30:0], main_spimaster3_spimachine3_sdi});
assign main_spimaster3_spimachine3_cnt_done = (main_spimaster3_spimachine3_cnt == 1'd0);
assign main_spimaster3_spimachine3_done = (main_spimaster3_spimachine3_cnt_done & (~main_spimaster3_spimachine3_do_extend));

// synthesis translate_off
reg dummy_d_84;
// synthesis translate_on
always @(*) begin
	main_spimaster3_spimachine3_clk_next <= 1'd0;
	main_spimaster3_spimachine3_cs_next <= 1'd0;
	main_spimaster3_spimachine3_idle <= 1'd0;
	main_spimaster3_spimachine3_readable <= 1'd0;
	main_spimaster3_spimachine3_writable <= 1'd0;
	main_spimaster3_spimachine3_load1 <= 1'd0;
	main_spimaster3_spimachine3_shift <= 1'd0;
	main_spimaster3_spimachine3_sample <= 1'd0;
	main_spimaster3_spimachine3_extend <= 1'd0;
	main_spimaster3_spimachine3_count <= 1'd0;
	builder_spimaster3_next_state <= 3'd0;
	builder_spimaster3_next_state <= builder_spimaster3_state;
	case (builder_spimaster3_state)
		1'd1: begin
			main_spimaster3_spimachine3_cs_next <= 1'd1;
			main_spimaster3_spimachine3_count <= 1'd1;
			main_spimaster3_spimachine3_extend <= 1'd1;
			main_spimaster3_spimachine3_clk_next <= 1'd1;
			if (main_spimaster3_spimachine3_done) begin
				builder_spimaster3_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster3_spimachine3_cs_next <= 1'd1;
			main_spimaster3_spimachine3_count <= 1'd1;
			main_spimaster3_spimachine3_clk_next <= (~main_spimaster3_spimachine3_clk_phase);
			if (main_spimaster3_spimachine3_done) begin
				main_spimaster3_spimachine3_sample <= 1'd1;
				builder_spimaster3_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster3_spimachine3_cs_next <= 1'd1;
			main_spimaster3_spimachine3_count <= 1'd1;
			main_spimaster3_spimachine3_extend <= 1'd1;
			main_spimaster3_spimachine3_clk_next <= main_spimaster3_spimachine3_clk_phase;
			if (main_spimaster3_spimachine3_done) begin
				if ((main_spimaster3_spimachine3_n == 1'd0)) begin
					main_spimaster3_spimachine3_readable <= 1'd1;
					main_spimaster3_spimachine3_writable <= 1'd1;
					if (main_spimaster3_spimachine3_end1) begin
						main_spimaster3_spimachine3_clk_next <= 1'd0;
						main_spimaster3_spimachine3_writable <= 1'd0;
						if (main_spimaster3_spimachine3_clk_phase) begin
							main_spimaster3_spimachine3_cs_next <= 1'd0;
							builder_spimaster3_next_state <= 3'd5;
						end else begin
							builder_spimaster3_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster3_spimachine3_load0) begin
							main_spimaster3_spimachine3_load1 <= 1'd1;
							builder_spimaster3_next_state <= 2'd2;
						end else begin
							main_spimaster3_spimachine3_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster3_spimachine3_shift <= 1'd1;
					builder_spimaster3_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster3_spimachine3_count <= 1'd1;
			if (main_spimaster3_spimachine3_done) begin
				builder_spimaster3_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster3_spimachine3_done) begin
				builder_spimaster3_next_state <= 1'd0;
			end else begin
				main_spimaster3_spimachine3_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster3_spimachine3_idle <= 1'd1;
			main_spimaster3_spimachine3_writable <= 1'd1;
			main_spimaster3_spimachine3_cs_next <= 1'd1;
			if (main_spimaster3_spimachine3_load0) begin
				main_spimaster3_spimachine3_count <= 1'd1;
				main_spimaster3_spimachine3_load1 <= 1'd1;
				if (main_spimaster3_spimachine3_clk_phase) begin
					builder_spimaster3_next_state <= 1'd1;
				end else begin
					main_spimaster3_spimachine3_extend <= 1'd1;
					builder_spimaster3_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_84 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster4_spimachine4_length = main_spimaster4_config_length;
assign main_spimaster4_spimachine4_end0 = main_spimaster4_config_end;
assign main_spimaster4_spimachine4_div = main_spimaster4_config_div;
assign main_spimaster4_spimachine4_clk_phase = main_spimaster4_config_clk_phase;
assign main_spimaster4_spimachine4_lsb_first = main_spimaster4_config_lsb_first;
assign main_spimaster4_interface_half_duplex = main_spimaster4_config_half_duplex;
assign main_spimaster4_interface_cs = main_spimaster4_config_cs;
assign main_spimaster4_interface_cs_polarity = {1{main_spimaster4_config_cs_polarity}};
assign main_spimaster4_interface_clk_polarity = main_spimaster4_config_clk_polarity;
assign main_spimaster4_interface_offline = main_spimaster4_config_offline;
assign main_spimaster4_interface_cs_next = main_spimaster4_spimachine4_cs_next;
assign main_spimaster4_interface_clk_next = main_spimaster4_spimachine4_clk_next;
assign main_spimaster4_interface_ce = main_spimaster4_spimachine4_ce;
assign main_spimaster4_interface_sample = main_spimaster4_spimachine4_sample;
assign main_spimaster4_spimachine4_sdi = main_spimaster4_interface_sdi;
assign main_spimaster4_interface_sdo = main_spimaster4_spimachine4_sdo;
assign main_spimaster4_spimachine4_load0 = ((main_spimaster4_ointerface4_stb & main_spimaster4_spimachine4_writable) & (~main_spimaster4_ointerface4_address));
assign main_spimaster4_spimachine4_pdo = main_spimaster4_ointerface4_data;
assign main_spimaster4_ointerface4_busy = (~main_spimaster4_spimachine4_writable);
assign main_spimaster4_iinterface4_stb = (main_spimaster4_spimachine4_readable & main_spimaster4_read);
assign main_spimaster4_iinterface4_data = main_spimaster4_spimachine4_pdi;
assign main_spimaster4_interface_miso_oe = 1'd0;
assign main_spimaster4_interface_mosi_o = main_spimaster4_interface_sdo;
assign main_spimaster4_interface_miso_o = main_spimaster4_interface_sdo;
assign main_spimaster4_interface_cs_oe = (~main_spimaster4_interface_offline);
assign main_spimaster4_interface_clk_oe = (~main_spimaster4_interface_offline);
assign main_spimaster4_interface_mosi_oe = (~(main_spimaster4_interface_offline | main_spimaster4_interface_half_duplex));

// synthesis translate_off
reg dummy_d_85;
// synthesis translate_on
always @(*) begin
	main_spimaster4_interface_sdi <= 1'd0;
	if ((main_spimaster4_interface_cs != 1'd0)) begin
		main_spimaster4_interface_sdi <= (main_spimaster4_interface_half_duplex ? main_spimaster4_interface_mosi_reg : main_spimaster4_interface_miso_reg);
	end
// synthesis translate_off
	dummy_d_85 <= dummy_s;
// synthesis translate_on
end
assign main_spimaster4_spimachine4_ce = (main_spimaster4_spimachine4_done & main_spimaster4_spimachine4_count);
assign main_spimaster4_spimachine4_pdi = (main_spimaster4_spimachine4_lsb_first ? {main_spimaster4_spimachine4_sdi, main_spimaster4_spimachine4_sr[31:1]} : {main_spimaster4_spimachine4_sr[30:0], main_spimaster4_spimachine4_sdi});
assign main_spimaster4_spimachine4_cnt_done = (main_spimaster4_spimachine4_cnt == 1'd0);
assign main_spimaster4_spimachine4_done = (main_spimaster4_spimachine4_cnt_done & (~main_spimaster4_spimachine4_do_extend));

// synthesis translate_off
reg dummy_d_86;
// synthesis translate_on
always @(*) begin
	main_spimaster4_spimachine4_clk_next <= 1'd0;
	main_spimaster4_spimachine4_cs_next <= 1'd0;
	main_spimaster4_spimachine4_idle <= 1'd0;
	main_spimaster4_spimachine4_readable <= 1'd0;
	main_spimaster4_spimachine4_writable <= 1'd0;
	main_spimaster4_spimachine4_load1 <= 1'd0;
	main_spimaster4_spimachine4_shift <= 1'd0;
	main_spimaster4_spimachine4_sample <= 1'd0;
	main_spimaster4_spimachine4_extend <= 1'd0;
	main_spimaster4_spimachine4_count <= 1'd0;
	builder_spimaster4_next_state <= 3'd0;
	builder_spimaster4_next_state <= builder_spimaster4_state;
	case (builder_spimaster4_state)
		1'd1: begin
			main_spimaster4_spimachine4_cs_next <= 1'd1;
			main_spimaster4_spimachine4_count <= 1'd1;
			main_spimaster4_spimachine4_extend <= 1'd1;
			main_spimaster4_spimachine4_clk_next <= 1'd1;
			if (main_spimaster4_spimachine4_done) begin
				builder_spimaster4_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_spimaster4_spimachine4_cs_next <= 1'd1;
			main_spimaster4_spimachine4_count <= 1'd1;
			main_spimaster4_spimachine4_clk_next <= (~main_spimaster4_spimachine4_clk_phase);
			if (main_spimaster4_spimachine4_done) begin
				main_spimaster4_spimachine4_sample <= 1'd1;
				builder_spimaster4_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_spimaster4_spimachine4_cs_next <= 1'd1;
			main_spimaster4_spimachine4_count <= 1'd1;
			main_spimaster4_spimachine4_extend <= 1'd1;
			main_spimaster4_spimachine4_clk_next <= main_spimaster4_spimachine4_clk_phase;
			if (main_spimaster4_spimachine4_done) begin
				if ((main_spimaster4_spimachine4_n == 1'd0)) begin
					main_spimaster4_spimachine4_readable <= 1'd1;
					main_spimaster4_spimachine4_writable <= 1'd1;
					if (main_spimaster4_spimachine4_end1) begin
						main_spimaster4_spimachine4_clk_next <= 1'd0;
						main_spimaster4_spimachine4_writable <= 1'd0;
						if (main_spimaster4_spimachine4_clk_phase) begin
							main_spimaster4_spimachine4_cs_next <= 1'd0;
							builder_spimaster4_next_state <= 3'd5;
						end else begin
							builder_spimaster4_next_state <= 3'd4;
						end
					end else begin
						if (main_spimaster4_spimachine4_load0) begin
							main_spimaster4_spimachine4_load1 <= 1'd1;
							builder_spimaster4_next_state <= 2'd2;
						end else begin
							main_spimaster4_spimachine4_count <= 1'd0;
						end
					end
				end else begin
					main_spimaster4_spimachine4_shift <= 1'd1;
					builder_spimaster4_next_state <= 2'd2;
				end
			end
		end
		3'd4: begin
			main_spimaster4_spimachine4_count <= 1'd1;
			if (main_spimaster4_spimachine4_done) begin
				builder_spimaster4_next_state <= 3'd5;
			end
		end
		3'd5: begin
			if (main_spimaster4_spimachine4_done) begin
				builder_spimaster4_next_state <= 1'd0;
			end else begin
				main_spimaster4_spimachine4_count <= 1'd1;
			end
		end
		default: begin
			main_spimaster4_spimachine4_idle <= 1'd1;
			main_spimaster4_spimachine4_writable <= 1'd1;
			main_spimaster4_spimachine4_cs_next <= 1'd1;
			if (main_spimaster4_spimachine4_load0) begin
				main_spimaster4_spimachine4_count <= 1'd1;
				main_spimaster4_spimachine4_load1 <= 1'd1;
				if (main_spimaster4_spimachine4_clk_phase) begin
					builder_spimaster4_next_state <= 1'd1;
				end else begin
					main_spimaster4_spimachine4_extend <= 1'd1;
					builder_spimaster4_next_state <= 2'd2;
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_86 <= dummy_s;
// synthesis translate_on
end
assign dds_rst = main_ad9914_gpio[0];
assign dds_sel_n = (~main_ad9914_gpio[11:1]);

// synthesis translate_off
reg dummy_d_87;
// synthesis translate_on
always @(*) begin
	main_ad9914_bus_dat_r <= 16'd0;
	if (main_ad9914_bus_r_gpio) begin
		main_ad9914_bus_dat_r <= main_ad9914_gpio;
	end else begin
		main_ad9914_bus_dat_r <= main_ad9914_dr;
	end
// synthesis translate_off
	dummy_d_87 <= dummy_s;
// synthesis translate_on
end
assign main_ad9914_read_timer_done = (main_ad9914_read_timer_count == 1'd0);
assign main_ad9914_hiz_timer_done = (main_ad9914_hiz_timer_count == 1'd0);

// synthesis translate_off
reg dummy_d_88;
// synthesis translate_on
always @(*) begin
	main_ad9914_bus_ack <= 1'd0;
	main_ad9914_hold_address <= 1'd0;
	main_ad9914_rx <= 1'd0;
	main_ad9914_gpio_load <= 1'd0;
	main_ad9914_bus_r_gpio <= 1'd0;
	main_ad9914_fud <= 1'd0;
	main_ad9914_wr <= 1'd0;
	main_ad9914_rd <= 1'd0;
	main_ad9914_read_timer_wait <= 1'd0;
	main_ad9914_hiz_timer_wait <= 1'd0;
	builder_ad9914_next_state <= 3'd0;
	builder_ad9914_next_state <= builder_ad9914_state;
	case (builder_ad9914_state)
		1'd1: begin
			main_ad9914_wr <= 1'd1;
			builder_ad9914_next_state <= 2'd2;
		end
		2'd2: begin
			main_ad9914_bus_ack <= 1'd1;
			builder_ad9914_next_state <= 1'd0;
		end
		2'd3: begin
			main_ad9914_rx <= 1'd1;
			main_ad9914_rd <= 1'd1;
			main_ad9914_read_timer_wait <= 1'd1;
			if (main_ad9914_read_timer_done) begin
				main_ad9914_bus_ack <= 1'd1;
				builder_ad9914_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_ad9914_rx <= 1'd1;
			main_ad9914_hold_address <= 1'd1;
			main_ad9914_hiz_timer_wait <= 1'd1;
			if (main_ad9914_hiz_timer_done) begin
				builder_ad9914_next_state <= 1'd0;
			end
		end
		3'd5: begin
			main_ad9914_fud <= 1'd1;
			main_ad9914_bus_ack <= 1'd1;
			builder_ad9914_next_state <= 1'd0;
		end
		3'd6: begin
			main_ad9914_bus_ack <= 1'd1;
			main_ad9914_bus_r_gpio <= 1'd1;
			if (main_ad9914_bus_we) begin
				main_ad9914_gpio_load <= 1'd1;
			end
			builder_ad9914_next_state <= 1'd0;
		end
		default: begin
			if ((main_ad9914_bus_cyc & main_ad9914_bus_stb)) begin
				if (main_ad9914_bus_adr[7]) begin
					if (main_ad9914_bus_adr[0]) begin
						builder_ad9914_next_state <= 3'd6;
					end else begin
						builder_ad9914_next_state <= 3'd5;
					end
				end else begin
					if (main_ad9914_bus_we) begin
						builder_ad9914_next_state <= 1'd1;
					end else begin
						builder_ad9914_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
// synthesis translate_off
	dummy_d_88 <= dummy_s;
// synthesis translate_on
end
assign main_ad9914_busy = main_ad9914_active;
assign main_ad9914_bus_cyc = main_ad9914_active;
assign main_ad9914_bus_stb = main_ad9914_active;
assign main_i = main_coarse_ts;
assign main_coarse_ts_sys = main_o;
assign main_full_ts = (main_coarse_ts <<< 2'd3);
assign main_full_ts_sys = (main_coarse_ts_sys <<< 2'd3);

// synthesis translate_off
reg dummy_d_89;
// synthesis translate_on
always @(*) begin
	main_value_sys <= 61'd0;
	main_value_sys[60] <= main_value_gray_sys[60];
	main_value_sys[59] <= (main_value_sys[60] ^ main_value_gray_sys[59]);
	main_value_sys[58] <= (main_value_sys[59] ^ main_value_gray_sys[58]);
	main_value_sys[57] <= (main_value_sys[58] ^ main_value_gray_sys[57]);
	main_value_sys[56] <= (main_value_sys[57] ^ main_value_gray_sys[56]);
	main_value_sys[55] <= (main_value_sys[56] ^ main_value_gray_sys[55]);
	main_value_sys[54] <= (main_value_sys[55] ^ main_value_gray_sys[54]);
	main_value_sys[53] <= (main_value_sys[54] ^ main_value_gray_sys[53]);
	main_value_sys[52] <= (main_value_sys[53] ^ main_value_gray_sys[52]);
	main_value_sys[51] <= (main_value_sys[52] ^ main_value_gray_sys[51]);
	main_value_sys[50] <= (main_value_sys[51] ^ main_value_gray_sys[50]);
	main_value_sys[49] <= (main_value_sys[50] ^ main_value_gray_sys[49]);
	main_value_sys[48] <= (main_value_sys[49] ^ main_value_gray_sys[48]);
	main_value_sys[47] <= (main_value_sys[48] ^ main_value_gray_sys[47]);
	main_value_sys[46] <= (main_value_sys[47] ^ main_value_gray_sys[46]);
	main_value_sys[45] <= (main_value_sys[46] ^ main_value_gray_sys[45]);
	main_value_sys[44] <= (main_value_sys[45] ^ main_value_gray_sys[44]);
	main_value_sys[43] <= (main_value_sys[44] ^ main_value_gray_sys[43]);
	main_value_sys[42] <= (main_value_sys[43] ^ main_value_gray_sys[42]);
	main_value_sys[41] <= (main_value_sys[42] ^ main_value_gray_sys[41]);
	main_value_sys[40] <= (main_value_sys[41] ^ main_value_gray_sys[40]);
	main_value_sys[39] <= (main_value_sys[40] ^ main_value_gray_sys[39]);
	main_value_sys[38] <= (main_value_sys[39] ^ main_value_gray_sys[38]);
	main_value_sys[37] <= (main_value_sys[38] ^ main_value_gray_sys[37]);
	main_value_sys[36] <= (main_value_sys[37] ^ main_value_gray_sys[36]);
	main_value_sys[35] <= (main_value_sys[36] ^ main_value_gray_sys[35]);
	main_value_sys[34] <= (main_value_sys[35] ^ main_value_gray_sys[34]);
	main_value_sys[33] <= (main_value_sys[34] ^ main_value_gray_sys[33]);
	main_value_sys[32] <= (main_value_sys[33] ^ main_value_gray_sys[32]);
	main_value_sys[31] <= (main_value_sys[32] ^ main_value_gray_sys[31]);
	main_value_sys[30] <= (main_value_sys[31] ^ main_value_gray_sys[30]);
	main_value_sys[29] <= (main_value_sys[30] ^ main_value_gray_sys[29]);
	main_value_sys[28] <= (main_value_sys[29] ^ main_value_gray_sys[28]);
	main_value_sys[27] <= (main_value_sys[28] ^ main_value_gray_sys[27]);
	main_value_sys[26] <= (main_value_sys[27] ^ main_value_gray_sys[26]);
	main_value_sys[25] <= (main_value_sys[26] ^ main_value_gray_sys[25]);
	main_value_sys[24] <= (main_value_sys[25] ^ main_value_gray_sys[24]);
	main_value_sys[23] <= (main_value_sys[24] ^ main_value_gray_sys[23]);
	main_value_sys[22] <= (main_value_sys[23] ^ main_value_gray_sys[22]);
	main_value_sys[21] <= (main_value_sys[22] ^ main_value_gray_sys[21]);
	main_value_sys[20] <= (main_value_sys[21] ^ main_value_gray_sys[20]);
	main_value_sys[19] <= (main_value_sys[20] ^ main_value_gray_sys[19]);
	main_value_sys[18] <= (main_value_sys[19] ^ main_value_gray_sys[18]);
	main_value_sys[17] <= (main_value_sys[18] ^ main_value_gray_sys[17]);
	main_value_sys[16] <= (main_value_sys[17] ^ main_value_gray_sys[16]);
	main_value_sys[15] <= (main_value_sys[16] ^ main_value_gray_sys[15]);
	main_value_sys[14] <= (main_value_sys[15] ^ main_value_gray_sys[14]);
	main_value_sys[13] <= (main_value_sys[14] ^ main_value_gray_sys[13]);
	main_value_sys[12] <= (main_value_sys[13] ^ main_value_gray_sys[12]);
	main_value_sys[11] <= (main_value_sys[12] ^ main_value_gray_sys[11]);
	main_value_sys[10] <= (main_value_sys[11] ^ main_value_gray_sys[10]);
	main_value_sys[9] <= (main_value_sys[10] ^ main_value_gray_sys[9]);
	main_value_sys[8] <= (main_value_sys[9] ^ main_value_gray_sys[8]);
	main_value_sys[7] <= (main_value_sys[8] ^ main_value_gray_sys[7]);
	main_value_sys[6] <= (main_value_sys[7] ^ main_value_gray_sys[6]);
	main_value_sys[5] <= (main_value_sys[6] ^ main_value_gray_sys[5]);
	main_value_sys[4] <= (main_value_sys[5] ^ main_value_gray_sys[4]);
	main_value_sys[3] <= (main_value_sys[4] ^ main_value_gray_sys[3]);
	main_value_sys[2] <= (main_value_sys[3] ^ main_value_gray_sys[2]);
	main_value_sys[1] <= (main_value_sys[2] ^ main_value_gray_sys[1]);
	main_value_sys[0] <= (main_value_sys[1] ^ main_value_gray_sys[0]);
// synthesis translate_off
	dummy_d_89 <= dummy_s;
// synthesis translate_on
end
assign rsys_clk = sys_clk;
assign rsys_rst = main_rtio_core_cmd_reset;
assign rio_clk = rtio_clk;
assign rio_phy_clk = rtio_clk;
assign main_rtio_core_outputs_gates_coarse_timestamp = main_coarse_ts;
assign main_rtio_core_async_error_w = {main_rtio_core_o_sequence_error, main_rtio_core_o_busy, main_rtio_core_o_collision};
assign main_rtio_core_o_collision_sync_i = main_rtio_core_outputs_collision;
assign main_rtio_core_o_collision_sync_data_i = main_rtio_core_outputs_collision_channel;
assign main_rtio_core_o_busy_sync_i = main_rtio_core_outputs_busy;
assign main_rtio_core_o_busy_sync_data_i = main_rtio_core_outputs_busy_channel;
assign main_rtio_core_outputs_record0_we = main_rtio_core_outputs_lanedistributor_record0_we;
assign main_rtio_core_outputs_lanedistributor_record0_writable = main_rtio_core_outputs_record0_writable;
assign main_rtio_core_outputs_record0_seqn0 = main_rtio_core_outputs_lanedistributor_record0_seqn;
assign main_rtio_core_outputs_record0_payload_channel0 = main_rtio_core_outputs_lanedistributor_record0_payload_channel;
assign main_rtio_core_outputs_record0_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record0_payload_timestamp;
assign main_rtio_core_outputs_record0_payload_address0 = main_rtio_core_outputs_lanedistributor_record0_payload_address;
assign main_rtio_core_outputs_record0_payload_data0 = main_rtio_core_outputs_lanedistributor_record0_payload_data;
assign main_rtio_core_outputs_record1_we = main_rtio_core_outputs_lanedistributor_record1_we;
assign main_rtio_core_outputs_lanedistributor_record1_writable = main_rtio_core_outputs_record1_writable;
assign main_rtio_core_outputs_record1_seqn0 = main_rtio_core_outputs_lanedistributor_record1_seqn;
assign main_rtio_core_outputs_record1_payload_channel0 = main_rtio_core_outputs_lanedistributor_record1_payload_channel;
assign main_rtio_core_outputs_record1_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record1_payload_timestamp;
assign main_rtio_core_outputs_record1_payload_address0 = main_rtio_core_outputs_lanedistributor_record1_payload_address;
assign main_rtio_core_outputs_record1_payload_data0 = main_rtio_core_outputs_lanedistributor_record1_payload_data;
assign main_rtio_core_outputs_record2_we = main_rtio_core_outputs_lanedistributor_record2_we;
assign main_rtio_core_outputs_lanedistributor_record2_writable = main_rtio_core_outputs_record2_writable;
assign main_rtio_core_outputs_record2_seqn0 = main_rtio_core_outputs_lanedistributor_record2_seqn;
assign main_rtio_core_outputs_record2_payload_channel0 = main_rtio_core_outputs_lanedistributor_record2_payload_channel;
assign main_rtio_core_outputs_record2_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record2_payload_timestamp;
assign main_rtio_core_outputs_record2_payload_address0 = main_rtio_core_outputs_lanedistributor_record2_payload_address;
assign main_rtio_core_outputs_record2_payload_data0 = main_rtio_core_outputs_lanedistributor_record2_payload_data;
assign main_rtio_core_outputs_record3_we = main_rtio_core_outputs_lanedistributor_record3_we;
assign main_rtio_core_outputs_lanedistributor_record3_writable = main_rtio_core_outputs_record3_writable;
assign main_rtio_core_outputs_record3_seqn0 = main_rtio_core_outputs_lanedistributor_record3_seqn;
assign main_rtio_core_outputs_record3_payload_channel0 = main_rtio_core_outputs_lanedistributor_record3_payload_channel;
assign main_rtio_core_outputs_record3_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record3_payload_timestamp;
assign main_rtio_core_outputs_record3_payload_address0 = main_rtio_core_outputs_lanedistributor_record3_payload_address;
assign main_rtio_core_outputs_record3_payload_data0 = main_rtio_core_outputs_lanedistributor_record3_payload_data;
assign main_rtio_core_outputs_record4_we = main_rtio_core_outputs_lanedistributor_record4_we;
assign main_rtio_core_outputs_lanedistributor_record4_writable = main_rtio_core_outputs_record4_writable;
assign main_rtio_core_outputs_record4_seqn0 = main_rtio_core_outputs_lanedistributor_record4_seqn;
assign main_rtio_core_outputs_record4_payload_channel0 = main_rtio_core_outputs_lanedistributor_record4_payload_channel;
assign main_rtio_core_outputs_record4_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record4_payload_timestamp;
assign main_rtio_core_outputs_record4_payload_address0 = main_rtio_core_outputs_lanedistributor_record4_payload_address;
assign main_rtio_core_outputs_record4_payload_data0 = main_rtio_core_outputs_lanedistributor_record4_payload_data;
assign main_rtio_core_outputs_record5_we = main_rtio_core_outputs_lanedistributor_record5_we;
assign main_rtio_core_outputs_lanedistributor_record5_writable = main_rtio_core_outputs_record5_writable;
assign main_rtio_core_outputs_record5_seqn0 = main_rtio_core_outputs_lanedistributor_record5_seqn;
assign main_rtio_core_outputs_record5_payload_channel0 = main_rtio_core_outputs_lanedistributor_record5_payload_channel;
assign main_rtio_core_outputs_record5_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record5_payload_timestamp;
assign main_rtio_core_outputs_record5_payload_address0 = main_rtio_core_outputs_lanedistributor_record5_payload_address;
assign main_rtio_core_outputs_record5_payload_data0 = main_rtio_core_outputs_lanedistributor_record5_payload_data;
assign main_rtio_core_outputs_record6_we = main_rtio_core_outputs_lanedistributor_record6_we;
assign main_rtio_core_outputs_lanedistributor_record6_writable = main_rtio_core_outputs_record6_writable;
assign main_rtio_core_outputs_record6_seqn0 = main_rtio_core_outputs_lanedistributor_record6_seqn;
assign main_rtio_core_outputs_record6_payload_channel0 = main_rtio_core_outputs_lanedistributor_record6_payload_channel;
assign main_rtio_core_outputs_record6_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record6_payload_timestamp;
assign main_rtio_core_outputs_record6_payload_address0 = main_rtio_core_outputs_lanedistributor_record6_payload_address;
assign main_rtio_core_outputs_record6_payload_data0 = main_rtio_core_outputs_lanedistributor_record6_payload_data;
assign main_rtio_core_outputs_record7_we = main_rtio_core_outputs_lanedistributor_record7_we;
assign main_rtio_core_outputs_lanedistributor_record7_writable = main_rtio_core_outputs_record7_writable;
assign main_rtio_core_outputs_record7_seqn0 = main_rtio_core_outputs_lanedistributor_record7_seqn;
assign main_rtio_core_outputs_record7_payload_channel0 = main_rtio_core_outputs_lanedistributor_record7_payload_channel;
assign main_rtio_core_outputs_record7_payload_timestamp0 = main_rtio_core_outputs_lanedistributor_record7_payload_timestamp;
assign main_rtio_core_outputs_record7_payload_address0 = main_rtio_core_outputs_lanedistributor_record7_payload_address;
assign main_rtio_core_outputs_record7_payload_data0 = main_rtio_core_outputs_lanedistributor_record7_payload_data;
assign main_rtio_core_outputs_record0_re = main_rtio_core_outputs_gates_record0_re;
assign main_rtio_core_outputs_gates_record0_readable = main_rtio_core_outputs_record0_readable;
assign main_rtio_core_outputs_gates_record0_seqn0 = main_rtio_core_outputs_record0_seqn1;
assign main_rtio_core_outputs_gates_record0_payload_channel0 = main_rtio_core_outputs_record0_payload_channel1;
assign main_rtio_core_outputs_gates_record0_payload_timestamp = main_rtio_core_outputs_record0_payload_timestamp1;
assign main_rtio_core_outputs_gates_record0_payload_address0 = main_rtio_core_outputs_record0_payload_address1;
assign main_rtio_core_outputs_gates_record0_payload_data0 = main_rtio_core_outputs_record0_payload_data1;
assign main_rtio_core_outputs_record1_re = main_rtio_core_outputs_gates_record1_re;
assign main_rtio_core_outputs_gates_record1_readable = main_rtio_core_outputs_record1_readable;
assign main_rtio_core_outputs_gates_record1_seqn0 = main_rtio_core_outputs_record1_seqn1;
assign main_rtio_core_outputs_gates_record1_payload_channel0 = main_rtio_core_outputs_record1_payload_channel1;
assign main_rtio_core_outputs_gates_record1_payload_timestamp = main_rtio_core_outputs_record1_payload_timestamp1;
assign main_rtio_core_outputs_gates_record1_payload_address0 = main_rtio_core_outputs_record1_payload_address1;
assign main_rtio_core_outputs_gates_record1_payload_data0 = main_rtio_core_outputs_record1_payload_data1;
assign main_rtio_core_outputs_record2_re = main_rtio_core_outputs_gates_record2_re;
assign main_rtio_core_outputs_gates_record2_readable = main_rtio_core_outputs_record2_readable;
assign main_rtio_core_outputs_gates_record2_seqn0 = main_rtio_core_outputs_record2_seqn1;
assign main_rtio_core_outputs_gates_record2_payload_channel0 = main_rtio_core_outputs_record2_payload_channel1;
assign main_rtio_core_outputs_gates_record2_payload_timestamp = main_rtio_core_outputs_record2_payload_timestamp1;
assign main_rtio_core_outputs_gates_record2_payload_address0 = main_rtio_core_outputs_record2_payload_address1;
assign main_rtio_core_outputs_gates_record2_payload_data0 = main_rtio_core_outputs_record2_payload_data1;
assign main_rtio_core_outputs_record3_re = main_rtio_core_outputs_gates_record3_re;
assign main_rtio_core_outputs_gates_record3_readable = main_rtio_core_outputs_record3_readable;
assign main_rtio_core_outputs_gates_record3_seqn0 = main_rtio_core_outputs_record3_seqn1;
assign main_rtio_core_outputs_gates_record3_payload_channel0 = main_rtio_core_outputs_record3_payload_channel1;
assign main_rtio_core_outputs_gates_record3_payload_timestamp = main_rtio_core_outputs_record3_payload_timestamp1;
assign main_rtio_core_outputs_gates_record3_payload_address0 = main_rtio_core_outputs_record3_payload_address1;
assign main_rtio_core_outputs_gates_record3_payload_data0 = main_rtio_core_outputs_record3_payload_data1;
assign main_rtio_core_outputs_record4_re = main_rtio_core_outputs_gates_record4_re;
assign main_rtio_core_outputs_gates_record4_readable = main_rtio_core_outputs_record4_readable;
assign main_rtio_core_outputs_gates_record4_seqn0 = main_rtio_core_outputs_record4_seqn1;
assign main_rtio_core_outputs_gates_record4_payload_channel0 = main_rtio_core_outputs_record4_payload_channel1;
assign main_rtio_core_outputs_gates_record4_payload_timestamp = main_rtio_core_outputs_record4_payload_timestamp1;
assign main_rtio_core_outputs_gates_record4_payload_address0 = main_rtio_core_outputs_record4_payload_address1;
assign main_rtio_core_outputs_gates_record4_payload_data0 = main_rtio_core_outputs_record4_payload_data1;
assign main_rtio_core_outputs_record5_re = main_rtio_core_outputs_gates_record5_re;
assign main_rtio_core_outputs_gates_record5_readable = main_rtio_core_outputs_record5_readable;
assign main_rtio_core_outputs_gates_record5_seqn0 = main_rtio_core_outputs_record5_seqn1;
assign main_rtio_core_outputs_gates_record5_payload_channel0 = main_rtio_core_outputs_record5_payload_channel1;
assign main_rtio_core_outputs_gates_record5_payload_timestamp = main_rtio_core_outputs_record5_payload_timestamp1;
assign main_rtio_core_outputs_gates_record5_payload_address0 = main_rtio_core_outputs_record5_payload_address1;
assign main_rtio_core_outputs_gates_record5_payload_data0 = main_rtio_core_outputs_record5_payload_data1;
assign main_rtio_core_outputs_record6_re = main_rtio_core_outputs_gates_record6_re;
assign main_rtio_core_outputs_gates_record6_readable = main_rtio_core_outputs_record6_readable;
assign main_rtio_core_outputs_gates_record6_seqn0 = main_rtio_core_outputs_record6_seqn1;
assign main_rtio_core_outputs_gates_record6_payload_channel0 = main_rtio_core_outputs_record6_payload_channel1;
assign main_rtio_core_outputs_gates_record6_payload_timestamp = main_rtio_core_outputs_record6_payload_timestamp1;
assign main_rtio_core_outputs_gates_record6_payload_address0 = main_rtio_core_outputs_record6_payload_address1;
assign main_rtio_core_outputs_gates_record6_payload_data0 = main_rtio_core_outputs_record6_payload_data1;
assign main_rtio_core_outputs_record7_re = main_rtio_core_outputs_gates_record7_re;
assign main_rtio_core_outputs_gates_record7_readable = main_rtio_core_outputs_record7_readable;
assign main_rtio_core_outputs_gates_record7_seqn0 = main_rtio_core_outputs_record7_seqn1;
assign main_rtio_core_outputs_gates_record7_payload_channel0 = main_rtio_core_outputs_record7_payload_channel1;
assign main_rtio_core_outputs_gates_record7_payload_timestamp = main_rtio_core_outputs_record7_payload_timestamp1;
assign main_rtio_core_outputs_gates_record7_payload_address0 = main_rtio_core_outputs_record7_payload_address1;
assign main_rtio_core_outputs_gates_record7_payload_data0 = main_rtio_core_outputs_record7_payload_data1;
assign main_rtio_core_outputs_record0_valid0 = main_rtio_core_outputs_gates_record0_valid;
assign main_rtio_core_outputs_record0_seqn2 = main_rtio_core_outputs_gates_record0_seqn1;
assign main_rtio_core_outputs_record0_replace_occured = main_rtio_core_outputs_gates_record0_replace_occured;
assign main_rtio_core_outputs_record0_nondata_replace_occured = main_rtio_core_outputs_gates_record0_nondata_replace_occured;
assign main_rtio_core_outputs_record0_payload_channel2 = main_rtio_core_outputs_gates_record0_payload_channel1;
assign main_rtio_core_outputs_record0_payload_fine_ts0 = main_rtio_core_outputs_gates_record0_payload_fine_ts;
assign main_rtio_core_outputs_record0_payload_address2 = main_rtio_core_outputs_gates_record0_payload_address1;
assign main_rtio_core_outputs_record0_payload_data2 = main_rtio_core_outputs_gates_record0_payload_data1;
assign main_rtio_core_outputs_record1_valid0 = main_rtio_core_outputs_gates_record1_valid;
assign main_rtio_core_outputs_record1_seqn2 = main_rtio_core_outputs_gates_record1_seqn1;
assign main_rtio_core_outputs_record1_replace_occured = main_rtio_core_outputs_gates_record1_replace_occured;
assign main_rtio_core_outputs_record1_nondata_replace_occured = main_rtio_core_outputs_gates_record1_nondata_replace_occured;
assign main_rtio_core_outputs_record1_payload_channel2 = main_rtio_core_outputs_gates_record1_payload_channel1;
assign main_rtio_core_outputs_record1_payload_fine_ts0 = main_rtio_core_outputs_gates_record1_payload_fine_ts;
assign main_rtio_core_outputs_record1_payload_address2 = main_rtio_core_outputs_gates_record1_payload_address1;
assign main_rtio_core_outputs_record1_payload_data2 = main_rtio_core_outputs_gates_record1_payload_data1;
assign main_rtio_core_outputs_record2_valid0 = main_rtio_core_outputs_gates_record2_valid;
assign main_rtio_core_outputs_record2_seqn2 = main_rtio_core_outputs_gates_record2_seqn1;
assign main_rtio_core_outputs_record2_replace_occured = main_rtio_core_outputs_gates_record2_replace_occured;
assign main_rtio_core_outputs_record2_nondata_replace_occured = main_rtio_core_outputs_gates_record2_nondata_replace_occured;
assign main_rtio_core_outputs_record2_payload_channel2 = main_rtio_core_outputs_gates_record2_payload_channel1;
assign main_rtio_core_outputs_record2_payload_fine_ts0 = main_rtio_core_outputs_gates_record2_payload_fine_ts;
assign main_rtio_core_outputs_record2_payload_address2 = main_rtio_core_outputs_gates_record2_payload_address1;
assign main_rtio_core_outputs_record2_payload_data2 = main_rtio_core_outputs_gates_record2_payload_data1;
assign main_rtio_core_outputs_record3_valid0 = main_rtio_core_outputs_gates_record3_valid;
assign main_rtio_core_outputs_record3_seqn2 = main_rtio_core_outputs_gates_record3_seqn1;
assign main_rtio_core_outputs_record3_replace_occured = main_rtio_core_outputs_gates_record3_replace_occured;
assign main_rtio_core_outputs_record3_nondata_replace_occured = main_rtio_core_outputs_gates_record3_nondata_replace_occured;
assign main_rtio_core_outputs_record3_payload_channel2 = main_rtio_core_outputs_gates_record3_payload_channel1;
assign main_rtio_core_outputs_record3_payload_fine_ts0 = main_rtio_core_outputs_gates_record3_payload_fine_ts;
assign main_rtio_core_outputs_record3_payload_address2 = main_rtio_core_outputs_gates_record3_payload_address1;
assign main_rtio_core_outputs_record3_payload_data2 = main_rtio_core_outputs_gates_record3_payload_data1;
assign main_rtio_core_outputs_record4_valid0 = main_rtio_core_outputs_gates_record4_valid;
assign main_rtio_core_outputs_record4_seqn2 = main_rtio_core_outputs_gates_record4_seqn1;
assign main_rtio_core_outputs_record4_replace_occured = main_rtio_core_outputs_gates_record4_replace_occured;
assign main_rtio_core_outputs_record4_nondata_replace_occured = main_rtio_core_outputs_gates_record4_nondata_replace_occured;
assign main_rtio_core_outputs_record4_payload_channel2 = main_rtio_core_outputs_gates_record4_payload_channel1;
assign main_rtio_core_outputs_record4_payload_fine_ts0 = main_rtio_core_outputs_gates_record4_payload_fine_ts;
assign main_rtio_core_outputs_record4_payload_address2 = main_rtio_core_outputs_gates_record4_payload_address1;
assign main_rtio_core_outputs_record4_payload_data2 = main_rtio_core_outputs_gates_record4_payload_data1;
assign main_rtio_core_outputs_record5_valid0 = main_rtio_core_outputs_gates_record5_valid;
assign main_rtio_core_outputs_record5_seqn2 = main_rtio_core_outputs_gates_record5_seqn1;
assign main_rtio_core_outputs_record5_replace_occured = main_rtio_core_outputs_gates_record5_replace_occured;
assign main_rtio_core_outputs_record5_nondata_replace_occured = main_rtio_core_outputs_gates_record5_nondata_replace_occured;
assign main_rtio_core_outputs_record5_payload_channel2 = main_rtio_core_outputs_gates_record5_payload_channel1;
assign main_rtio_core_outputs_record5_payload_fine_ts0 = main_rtio_core_outputs_gates_record5_payload_fine_ts;
assign main_rtio_core_outputs_record5_payload_address2 = main_rtio_core_outputs_gates_record5_payload_address1;
assign main_rtio_core_outputs_record5_payload_data2 = main_rtio_core_outputs_gates_record5_payload_data1;
assign main_rtio_core_outputs_record6_valid0 = main_rtio_core_outputs_gates_record6_valid;
assign main_rtio_core_outputs_record6_seqn2 = main_rtio_core_outputs_gates_record6_seqn1;
assign main_rtio_core_outputs_record6_replace_occured = main_rtio_core_outputs_gates_record6_replace_occured;
assign main_rtio_core_outputs_record6_nondata_replace_occured = main_rtio_core_outputs_gates_record6_nondata_replace_occured;
assign main_rtio_core_outputs_record6_payload_channel2 = main_rtio_core_outputs_gates_record6_payload_channel1;
assign main_rtio_core_outputs_record6_payload_fine_ts0 = main_rtio_core_outputs_gates_record6_payload_fine_ts;
assign main_rtio_core_outputs_record6_payload_address2 = main_rtio_core_outputs_gates_record6_payload_address1;
assign main_rtio_core_outputs_record6_payload_data2 = main_rtio_core_outputs_gates_record6_payload_data1;
assign main_rtio_core_outputs_record7_valid0 = main_rtio_core_outputs_gates_record7_valid;
assign main_rtio_core_outputs_record7_seqn2 = main_rtio_core_outputs_gates_record7_seqn1;
assign main_rtio_core_outputs_record7_replace_occured = main_rtio_core_outputs_gates_record7_replace_occured;
assign main_rtio_core_outputs_record7_nondata_replace_occured = main_rtio_core_outputs_gates_record7_nondata_replace_occured;
assign main_rtio_core_outputs_record7_payload_channel2 = main_rtio_core_outputs_gates_record7_payload_channel1;
assign main_rtio_core_outputs_record7_payload_fine_ts0 = main_rtio_core_outputs_gates_record7_payload_fine_ts;
assign main_rtio_core_outputs_record7_payload_address2 = main_rtio_core_outputs_gates_record7_payload_address1;
assign main_rtio_core_outputs_record7_payload_data2 = main_rtio_core_outputs_gates_record7_payload_data1;
assign main_rtio_core_cri_o_status = {main_rtio_core_outputs_lanedistributor_o_status_underflow, main_rtio_core_outputs_lanedistributor_o_status_wait};
assign main_rtio_core_outputs_lanedistributor_record0_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record0_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record0_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record0_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record1_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record1_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record1_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record1_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record2_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record2_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record2_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record2_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record3_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record3_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record3_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record3_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record4_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record4_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record4_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record4_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record5_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record5_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record5_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record5_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record6_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record6_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record6_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record6_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_record7_seqn = main_rtio_core_outputs_lanedistributor_seqn;
assign main_rtio_core_outputs_lanedistributor_record7_payload_channel = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_record7_payload_address = main_rtio_core_cri_o_address;
assign main_rtio_core_outputs_lanedistributor_record7_payload_data = main_rtio_core_cri_o_data;
assign main_rtio_core_outputs_lanedistributor_coarse_timestamp = main_rtio_core_cri_o_timestamp[63:3];
assign main_rtio_core_outputs_lanedistributor_current_lane_plus_one = (main_rtio_core_outputs_lanedistributor_current_lane + 1'd1);
assign main_rtio_core_outputs_lanedistributor_adr = main_rtio_core_cri_chan_sel[15:0];
assign main_rtio_core_outputs_lanedistributor_compensation = main_rtio_core_outputs_lanedistributor_dat_r;
assign main_rtio_core_outputs_lanedistributor_timestamp_above_min = ((main_rtio_core_outputs_lanedistributor_min_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min = ((main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min = ((main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));
assign main_rtio_core_outputs_lanedistributor_timestamp_above_last = ((main_rtio_core_outputs_lanedistributor_last_minus_timestamp - main_rtio_core_outputs_lanedistributor_compensation) < $signed({1'd0, 1'd0}));

// synthesis translate_off
reg dummy_d_90;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	main_rtio_core_outputs_lanedistributor_use_lanen <= 3'd0;
	if ((main_rtio_core_outputs_lanedistributor_force_laneB | (~main_rtio_core_outputs_lanedistributor_timestamp_above_last))) begin
		main_rtio_core_outputs_lanedistributor_use_lanen <= main_rtio_core_outputs_lanedistributor_current_lane_plus_one;
		main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd1;
	end else begin
		main_rtio_core_outputs_lanedistributor_use_lanen <= main_rtio_core_outputs_lanedistributor_current_lane;
		main_rtio_core_outputs_lanedistributor_use_laneB <= 1'd0;
	end
// synthesis translate_off
	dummy_d_90 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min = (main_rtio_core_outputs_lanedistributor_use_laneB ? main_rtio_core_outputs_lanedistributor_timestamp_above_laneB_min : main_rtio_core_outputs_lanedistributor_timestamp_above_laneA_min);

// synthesis translate_off
reg dummy_d_91;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_do_write <= 1'd0;
	main_rtio_core_outputs_lanedistributor_do_underflow <= 1'd0;
	main_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd0;
	if (((~main_rtio_core_outputs_lanedistributor_quash) & (main_rtio_core_cri_cmd == 1'd1))) begin
		if (main_rtio_core_outputs_lanedistributor_timestamp_above_min) begin
			if (main_rtio_core_outputs_lanedistributor_timestamp_above_lane_min) begin
				main_rtio_core_outputs_lanedistributor_do_write <= 1'd1;
			end else begin
				main_rtio_core_outputs_lanedistributor_do_sequence_error <= 1'd1;
			end
		end else begin
			main_rtio_core_outputs_lanedistributor_do_underflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_91 <= dummy_s;
// synthesis translate_on
end
assign builder_comb_lhs_array_muxed = main_rtio_core_outputs_lanedistributor_do_write;

// synthesis translate_off
reg dummy_d_92;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record0_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record1_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record2_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record3_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record4_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record5_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record6_we <= 1'd0;
	main_rtio_core_outputs_lanedistributor_record7_we <= 1'd0;
	case (main_rtio_core_outputs_lanedistributor_use_lanen)
		1'd0: begin
			main_rtio_core_outputs_lanedistributor_record0_we <= builder_comb_lhs_array_muxed;
		end
		1'd1: begin
			main_rtio_core_outputs_lanedistributor_record1_we <= builder_comb_lhs_array_muxed;
		end
		2'd2: begin
			main_rtio_core_outputs_lanedistributor_record2_we <= builder_comb_lhs_array_muxed;
		end
		2'd3: begin
			main_rtio_core_outputs_lanedistributor_record3_we <= builder_comb_lhs_array_muxed;
		end
		3'd4: begin
			main_rtio_core_outputs_lanedistributor_record4_we <= builder_comb_lhs_array_muxed;
		end
		3'd5: begin
			main_rtio_core_outputs_lanedistributor_record5_we <= builder_comb_lhs_array_muxed;
		end
		3'd6: begin
			main_rtio_core_outputs_lanedistributor_record6_we <= builder_comb_lhs_array_muxed;
		end
		default: begin
			main_rtio_core_outputs_lanedistributor_record7_we <= builder_comb_lhs_array_muxed;
		end
	endcase
// synthesis translate_off
	dummy_d_92 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_compensated_timestamp = ($signed({1'd0, main_rtio_core_cri_o_timestamp}) + (main_rtio_core_outputs_lanedistributor_compensation <<< 2'd3));

// synthesis translate_off
reg dummy_d_93;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record0_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_93 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_94;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record1_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_94 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_95;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record2_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_95 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_96;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record3_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_96 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_97;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record4_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_97 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_98;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record5_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_98 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_99;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record6_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_99 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_100;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= 64'd0;
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= main_rtio_core_cri_o_timestamp;
	main_rtio_core_outputs_lanedistributor_record7_payload_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp;
// synthesis translate_off
	dummy_d_100 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_lanedistributor_current_lane_writable = builder_comb_rhs_array_muxed8;
assign main_rtio_core_outputs_lanedistributor_o_status_wait = (~main_rtio_core_outputs_lanedistributor_current_lane_writable);
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din = {{main_rtio_core_outputs_record0_payload_data0, main_rtio_core_outputs_record0_payload_address0, main_rtio_core_outputs_record0_payload_timestamp0, main_rtio_core_outputs_record0_payload_channel0}, main_rtio_core_outputs_record0_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we = main_rtio_core_outputs_record0_we;
assign main_rtio_core_outputs_record0_writable = main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable;
assign {{main_rtio_core_outputs_record0_payload_data1, main_rtio_core_outputs_record0_payload_address1, main_rtio_core_outputs_record0_payload_timestamp1, main_rtio_core_outputs_record0_payload_channel1}, main_rtio_core_outputs_record0_seqn1} = main_rtio_core_outputs_asyncfifobuffered0_dout;
assign main_rtio_core_outputs_record0_readable = main_rtio_core_outputs_asyncfifobuffered0_readable;
assign main_rtio_core_outputs_asyncfifobuffered0_re = main_rtio_core_outputs_record0_re;
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din = {{main_rtio_core_outputs_record1_payload_data0, main_rtio_core_outputs_record1_payload_address0, main_rtio_core_outputs_record1_payload_timestamp0, main_rtio_core_outputs_record1_payload_channel0}, main_rtio_core_outputs_record1_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we = main_rtio_core_outputs_record1_we;
assign main_rtio_core_outputs_record1_writable = main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable;
assign {{main_rtio_core_outputs_record1_payload_data1, main_rtio_core_outputs_record1_payload_address1, main_rtio_core_outputs_record1_payload_timestamp1, main_rtio_core_outputs_record1_payload_channel1}, main_rtio_core_outputs_record1_seqn1} = main_rtio_core_outputs_asyncfifobuffered1_dout;
assign main_rtio_core_outputs_record1_readable = main_rtio_core_outputs_asyncfifobuffered1_readable;
assign main_rtio_core_outputs_asyncfifobuffered1_re = main_rtio_core_outputs_record1_re;
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din = {{main_rtio_core_outputs_record2_payload_data0, main_rtio_core_outputs_record2_payload_address0, main_rtio_core_outputs_record2_payload_timestamp0, main_rtio_core_outputs_record2_payload_channel0}, main_rtio_core_outputs_record2_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we = main_rtio_core_outputs_record2_we;
assign main_rtio_core_outputs_record2_writable = main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable;
assign {{main_rtio_core_outputs_record2_payload_data1, main_rtio_core_outputs_record2_payload_address1, main_rtio_core_outputs_record2_payload_timestamp1, main_rtio_core_outputs_record2_payload_channel1}, main_rtio_core_outputs_record2_seqn1} = main_rtio_core_outputs_asyncfifobuffered2_dout;
assign main_rtio_core_outputs_record2_readable = main_rtio_core_outputs_asyncfifobuffered2_readable;
assign main_rtio_core_outputs_asyncfifobuffered2_re = main_rtio_core_outputs_record2_re;
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din = {{main_rtio_core_outputs_record3_payload_data0, main_rtio_core_outputs_record3_payload_address0, main_rtio_core_outputs_record3_payload_timestamp0, main_rtio_core_outputs_record3_payload_channel0}, main_rtio_core_outputs_record3_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we = main_rtio_core_outputs_record3_we;
assign main_rtio_core_outputs_record3_writable = main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable;
assign {{main_rtio_core_outputs_record3_payload_data1, main_rtio_core_outputs_record3_payload_address1, main_rtio_core_outputs_record3_payload_timestamp1, main_rtio_core_outputs_record3_payload_channel1}, main_rtio_core_outputs_record3_seqn1} = main_rtio_core_outputs_asyncfifobuffered3_dout;
assign main_rtio_core_outputs_record3_readable = main_rtio_core_outputs_asyncfifobuffered3_readable;
assign main_rtio_core_outputs_asyncfifobuffered3_re = main_rtio_core_outputs_record3_re;
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din = {{main_rtio_core_outputs_record4_payload_data0, main_rtio_core_outputs_record4_payload_address0, main_rtio_core_outputs_record4_payload_timestamp0, main_rtio_core_outputs_record4_payload_channel0}, main_rtio_core_outputs_record4_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we = main_rtio_core_outputs_record4_we;
assign main_rtio_core_outputs_record4_writable = main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable;
assign {{main_rtio_core_outputs_record4_payload_data1, main_rtio_core_outputs_record4_payload_address1, main_rtio_core_outputs_record4_payload_timestamp1, main_rtio_core_outputs_record4_payload_channel1}, main_rtio_core_outputs_record4_seqn1} = main_rtio_core_outputs_asyncfifobuffered4_dout;
assign main_rtio_core_outputs_record4_readable = main_rtio_core_outputs_asyncfifobuffered4_readable;
assign main_rtio_core_outputs_asyncfifobuffered4_re = main_rtio_core_outputs_record4_re;
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din = {{main_rtio_core_outputs_record5_payload_data0, main_rtio_core_outputs_record5_payload_address0, main_rtio_core_outputs_record5_payload_timestamp0, main_rtio_core_outputs_record5_payload_channel0}, main_rtio_core_outputs_record5_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we = main_rtio_core_outputs_record5_we;
assign main_rtio_core_outputs_record5_writable = main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable;
assign {{main_rtio_core_outputs_record5_payload_data1, main_rtio_core_outputs_record5_payload_address1, main_rtio_core_outputs_record5_payload_timestamp1, main_rtio_core_outputs_record5_payload_channel1}, main_rtio_core_outputs_record5_seqn1} = main_rtio_core_outputs_asyncfifobuffered5_dout;
assign main_rtio_core_outputs_record5_readable = main_rtio_core_outputs_asyncfifobuffered5_readable;
assign main_rtio_core_outputs_asyncfifobuffered5_re = main_rtio_core_outputs_record5_re;
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din = {{main_rtio_core_outputs_record6_payload_data0, main_rtio_core_outputs_record6_payload_address0, main_rtio_core_outputs_record6_payload_timestamp0, main_rtio_core_outputs_record6_payload_channel0}, main_rtio_core_outputs_record6_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we = main_rtio_core_outputs_record6_we;
assign main_rtio_core_outputs_record6_writable = main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable;
assign {{main_rtio_core_outputs_record6_payload_data1, main_rtio_core_outputs_record6_payload_address1, main_rtio_core_outputs_record6_payload_timestamp1, main_rtio_core_outputs_record6_payload_channel1}, main_rtio_core_outputs_record6_seqn1} = main_rtio_core_outputs_asyncfifobuffered6_dout;
assign main_rtio_core_outputs_record6_readable = main_rtio_core_outputs_asyncfifobuffered6_readable;
assign main_rtio_core_outputs_asyncfifobuffered6_re = main_rtio_core_outputs_record6_re;
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din = {{main_rtio_core_outputs_record7_payload_data0, main_rtio_core_outputs_record7_payload_address0, main_rtio_core_outputs_record7_payload_timestamp0, main_rtio_core_outputs_record7_payload_channel0}, main_rtio_core_outputs_record7_seqn0};
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we = main_rtio_core_outputs_record7_we;
assign main_rtio_core_outputs_record7_writable = main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable;
assign {{main_rtio_core_outputs_record7_payload_data1, main_rtio_core_outputs_record7_payload_address1, main_rtio_core_outputs_record7_payload_timestamp1, main_rtio_core_outputs_record7_payload_channel1}, main_rtio_core_outputs_record7_seqn1} = main_rtio_core_outputs_asyncfifobuffered7_dout;
assign main_rtio_core_outputs_record7_readable = main_rtio_core_outputs_asyncfifobuffered7_readable;
assign main_rtio_core_outputs_asyncfifobuffered7_re = main_rtio_core_outputs_record7_re;
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re = (main_rtio_core_outputs_asyncfifobuffered0_re | (~main_rtio_core_outputs_asyncfifobuffered0_readable));
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce = (main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable & main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_we);
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce = (main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable & main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_re);
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_writable = (((main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[7] == main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[6] == main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q[5:0] != main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable = (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q != main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_adr = main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_din;
assign main_rtio_core_outputs_asyncfifobuffered0_wrport_we = main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce;
assign main_rtio_core_outputs_asyncfifobuffered0_rdport_adr = main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout = main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_101;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_ce) begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_101 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next = (main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_102;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_ce) begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_102 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next = (main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re = (main_rtio_core_outputs_asyncfifobuffered1_re | (~main_rtio_core_outputs_asyncfifobuffered1_readable));
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce = (main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable & main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_we);
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce = (main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable & main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_re);
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_writable = (((main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[7] == main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[6] == main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q[5:0] != main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable = (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q != main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_adr = main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_din;
assign main_rtio_core_outputs_asyncfifobuffered1_wrport_we = main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce;
assign main_rtio_core_outputs_asyncfifobuffered1_rdport_adr = main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout = main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_103;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_ce) begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_103 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next = (main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_104;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_ce) begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_104 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next = (main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re = (main_rtio_core_outputs_asyncfifobuffered2_re | (~main_rtio_core_outputs_asyncfifobuffered2_readable));
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce = (main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable & main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_we);
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce = (main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable & main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_re);
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_writable = (((main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[7] == main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[6] == main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q[5:0] != main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable = (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q != main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_adr = main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_din;
assign main_rtio_core_outputs_asyncfifobuffered2_wrport_we = main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce;
assign main_rtio_core_outputs_asyncfifobuffered2_rdport_adr = main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout = main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_105;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_ce) begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_105 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next = (main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_106;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_ce) begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_106 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next = (main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re = (main_rtio_core_outputs_asyncfifobuffered3_re | (~main_rtio_core_outputs_asyncfifobuffered3_readable));
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce = (main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable & main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_we);
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce = (main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable & main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_re);
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_writable = (((main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[7] == main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[6] == main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q[5:0] != main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable = (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q != main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_adr = main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_din;
assign main_rtio_core_outputs_asyncfifobuffered3_wrport_we = main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce;
assign main_rtio_core_outputs_asyncfifobuffered3_rdport_adr = main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout = main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_107;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_ce) begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_107 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next = (main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_108;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_ce) begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_108 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next = (main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re = (main_rtio_core_outputs_asyncfifobuffered4_re | (~main_rtio_core_outputs_asyncfifobuffered4_readable));
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce = (main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable & main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_we);
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce = (main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable & main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_re);
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_writable = (((main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[7] == main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[6] == main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q[5:0] != main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable = (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q != main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_adr = main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_din;
assign main_rtio_core_outputs_asyncfifobuffered4_wrport_we = main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce;
assign main_rtio_core_outputs_asyncfifobuffered4_rdport_adr = main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout = main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_109;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_ce) begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_109 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next = (main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_110;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_ce) begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_110 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next = (main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re = (main_rtio_core_outputs_asyncfifobuffered5_re | (~main_rtio_core_outputs_asyncfifobuffered5_readable));
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce = (main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable & main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_we);
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce = (main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable & main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_re);
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_writable = (((main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[7] == main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[6] == main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q[5:0] != main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable = (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q != main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_adr = main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_din;
assign main_rtio_core_outputs_asyncfifobuffered5_wrport_we = main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce;
assign main_rtio_core_outputs_asyncfifobuffered5_rdport_adr = main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout = main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_111;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_ce) begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_111 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next = (main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_112;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_ce) begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_112 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next = (main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re = (main_rtio_core_outputs_asyncfifobuffered6_re | (~main_rtio_core_outputs_asyncfifobuffered6_readable));
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce = (main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable & main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_we);
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce = (main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable & main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_re);
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_writable = (((main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[7] == main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[6] == main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q[5:0] != main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable = (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q != main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_adr = main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_din;
assign main_rtio_core_outputs_asyncfifobuffered6_wrport_we = main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce;
assign main_rtio_core_outputs_asyncfifobuffered6_rdport_adr = main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout = main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_113;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_ce) begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_113 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next = (main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_114;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_ce) begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_114 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next = (main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary[7:1]);
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re = (main_rtio_core_outputs_asyncfifobuffered7_re | (~main_rtio_core_outputs_asyncfifobuffered7_readable));
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce = (main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable & main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_we);
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce = (main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable & main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_re);
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_writable = (((main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[7] == main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[7]) | (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[6] == main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[6])) | (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q[5:0] != main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain[5:0]));
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable = (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q != main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain);
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_adr = main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w = main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_din;
assign main_rtio_core_outputs_asyncfifobuffered7_wrport_we = main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce;
assign main_rtio_core_outputs_asyncfifobuffered7_rdport_adr = main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[6:0];
assign main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout = main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r;

// synthesis translate_off
reg dummy_d_115;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_ce) begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary;
	end
// synthesis translate_off
	dummy_d_115 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next = (main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_116;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= 8'd0;
	if (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_ce) begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary + 1'd1);
	end else begin
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary;
	end
// synthesis translate_off
	dummy_d_116 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next = (main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary ^ main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary[7:1]);
assign main_rtio_core_outputs_gates_record0_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record0_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record0_re = (main_rtio_core_outputs_gates_record0_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record1_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record1_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record1_re = (main_rtio_core_outputs_gates_record1_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record2_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record2_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record2_re = (main_rtio_core_outputs_gates_record2_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record3_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record3_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record3_re = (main_rtio_core_outputs_gates_record3_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record4_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record4_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record4_re = (main_rtio_core_outputs_gates_record4_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record5_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record5_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record5_re = (main_rtio_core_outputs_gates_record5_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record6_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record6_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record6_re = (main_rtio_core_outputs_gates_record6_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_gates_record7_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record7_nondata_replace_occured = 1'd0;
assign main_rtio_core_outputs_gates_record7_re = (main_rtio_core_outputs_gates_record7_payload_timestamp[63:3] == main_rtio_core_outputs_gates_coarse_timestamp);
assign main_rtio_core_outputs_memory0_adr = main_rtio_core_outputs_record40_rec_payload_channel;
assign main_rtio_core_outputs_record0_collision = (main_rtio_core_outputs_replace_occured_r0 & ((~main_rtio_core_outputs_memory0_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r0));
assign main_rtio_core_outputs_memory1_adr = main_rtio_core_outputs_record41_rec_payload_channel;
assign main_rtio_core_outputs_record1_collision = (main_rtio_core_outputs_replace_occured_r1 & ((~main_rtio_core_outputs_memory1_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r1));
assign main_rtio_core_outputs_memory2_adr = main_rtio_core_outputs_record42_rec_payload_channel;
assign main_rtio_core_outputs_record2_collision = (main_rtio_core_outputs_replace_occured_r2 & ((~main_rtio_core_outputs_memory2_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r2));
assign main_rtio_core_outputs_memory3_adr = main_rtio_core_outputs_record43_rec_payload_channel;
assign main_rtio_core_outputs_record3_collision = (main_rtio_core_outputs_replace_occured_r3 & ((~main_rtio_core_outputs_memory3_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r3));
assign main_rtio_core_outputs_memory4_adr = main_rtio_core_outputs_record44_rec_payload_channel;
assign main_rtio_core_outputs_record4_collision = (main_rtio_core_outputs_replace_occured_r4 & ((~main_rtio_core_outputs_memory4_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r4));
assign main_rtio_core_outputs_memory5_adr = main_rtio_core_outputs_record45_rec_payload_channel;
assign main_rtio_core_outputs_record5_collision = (main_rtio_core_outputs_replace_occured_r5 & ((~main_rtio_core_outputs_memory5_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r5));
assign main_rtio_core_outputs_memory6_adr = main_rtio_core_outputs_record46_rec_payload_channel;
assign main_rtio_core_outputs_record6_collision = (main_rtio_core_outputs_replace_occured_r6 & ((~main_rtio_core_outputs_memory6_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r6));
assign main_rtio_core_outputs_memory7_adr = main_rtio_core_outputs_record47_rec_payload_channel;
assign main_rtio_core_outputs_record7_collision = (main_rtio_core_outputs_replace_occured_r7 & ((~main_rtio_core_outputs_memory7_dat_r) | main_rtio_core_outputs_nondata_replace_occured_r7));
assign main_rtio_core_outputs_selected0 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected1 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected2 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected3 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected4 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected5 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected6 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected7 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 1'd0));
assign main_rtio_core_outputs_selected8 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected9 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected10 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected11 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected12 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected13 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected14 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected15 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 1'd1));
assign main_rtio_core_outputs_selected16 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected17 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected18 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected19 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected20 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected21 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected22 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected23 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 2'd2));
assign main_rtio_core_outputs_selected24 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected25 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected26 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected27 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected28 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected29 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected30 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected31 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 2'd3));
assign main_rtio_core_outputs_selected32 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected33 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected34 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected35 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected36 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected37 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected38 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected39 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd4));
assign main_rtio_core_outputs_selected40 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected41 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected42 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected43 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected44 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected45 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected46 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected47 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd5));
assign main_rtio_core_outputs_selected48 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected49 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected50 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected51 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected52 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected53 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected54 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected55 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd6));
assign main_rtio_core_outputs_selected56 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected57 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected58 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected59 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected60 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected61 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected62 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected63 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 3'd7));
assign main_rtio_core_outputs_selected64 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected65 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected66 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected67 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected68 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected69 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected70 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected71 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd8));
assign main_rtio_core_outputs_selected72 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected73 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected74 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected75 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected76 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected77 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected78 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected79 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd9));
assign main_rtio_core_outputs_selected80 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected81 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected82 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected83 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected84 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected85 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected86 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected87 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd10));
assign main_rtio_core_outputs_selected88 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected89 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected90 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected91 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected92 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected93 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected94 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected95 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd11));
assign main_rtio_core_outputs_selected96 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected97 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected98 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected99 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected100 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected101 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected102 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected103 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd12));
assign main_rtio_core_outputs_selected104 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected105 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected106 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected107 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected108 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected109 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected110 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected111 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd13));
assign main_rtio_core_outputs_selected112 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected113 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected114 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected115 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected116 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected117 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected118 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected119 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd14));
assign main_rtio_core_outputs_selected120 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected121 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected122 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected123 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected124 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected125 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected126 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected127 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 4'd15));
assign main_rtio_core_outputs_selected128 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected129 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected130 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected131 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected132 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected133 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected134 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected135 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd16));
assign main_rtio_core_outputs_selected136 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected137 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected138 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected139 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected140 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected141 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected142 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected143 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd17));
assign main_rtio_core_outputs_selected144 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected145 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected146 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected147 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected148 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected149 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected150 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected151 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd18));
assign main_rtio_core_outputs_selected152 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected153 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected154 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected155 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected156 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected157 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected158 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected159 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd19));
assign main_rtio_core_outputs_selected160 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected161 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected162 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected163 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected164 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected165 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected166 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected167 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd20));
assign main_rtio_core_outputs_selected168 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected169 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected170 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected171 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected172 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected173 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected174 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected175 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd21));
assign main_rtio_core_outputs_selected176 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected177 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected178 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected179 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected180 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected181 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected182 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected183 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd22));
assign main_rtio_core_outputs_selected184 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected185 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected186 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected187 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected188 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected189 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected190 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected191 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd23));
assign main_rtio_core_outputs_selected192 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected193 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected194 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected195 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected196 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected197 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected198 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected199 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd24));
assign main_rtio_core_outputs_selected200 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected201 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected202 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected203 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected204 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected205 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected206 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected207 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd25));
assign main_rtio_core_outputs_selected208 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected209 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected210 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected211 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected212 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected213 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected214 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected215 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd26));
assign main_rtio_core_outputs_selected216 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected217 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected218 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected219 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected220 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected221 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected222 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected223 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd27));
assign main_rtio_core_outputs_selected224 = ((main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision)) & (main_rtio_core_outputs_record0_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected225 = ((main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision)) & (main_rtio_core_outputs_record1_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected226 = ((main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision)) & (main_rtio_core_outputs_record2_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected227 = ((main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision)) & (main_rtio_core_outputs_record3_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected228 = ((main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision)) & (main_rtio_core_outputs_record4_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected229 = ((main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision)) & (main_rtio_core_outputs_record5_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected230 = ((main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision)) & (main_rtio_core_outputs_record6_payload_channel3 == 5'd28));
assign main_rtio_core_outputs_selected231 = ((main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision)) & (main_rtio_core_outputs_record7_payload_channel3 == 5'd28));

// synthesis translate_off
reg dummy_d_117;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference0 <= 1'd0;
	if ((main_rtio_core_outputs_record0_payload_channel2 != main_rtio_core_outputs_record1_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_payload_fine_ts0 != main_rtio_core_outputs_record1_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_payload_address2 != main_rtio_core_outputs_record1_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference0 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_117 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_118;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference1 <= 1'd0;
	if ((main_rtio_core_outputs_record2_payload_channel2 != main_rtio_core_outputs_record3_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record2_payload_fine_ts0 != main_rtio_core_outputs_record3_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record2_payload_address2 != main_rtio_core_outputs_record3_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference1 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_118 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_119;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference2 <= 1'd0;
	if ((main_rtio_core_outputs_record4_payload_channel2 != main_rtio_core_outputs_record5_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_payload_fine_ts0 != main_rtio_core_outputs_record5_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_payload_address2 != main_rtio_core_outputs_record5_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference2 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_119 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_120;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference3 <= 1'd0;
	if ((main_rtio_core_outputs_record6_payload_channel2 != main_rtio_core_outputs_record7_payload_channel2)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record6_payload_fine_ts0 != main_rtio_core_outputs_record7_payload_fine_ts0)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record6_payload_address2 != main_rtio_core_outputs_record7_payload_address2)) begin
		main_rtio_core_outputs_nondata_difference3 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_120 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_121;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference4 <= 1'd0;
	if ((main_rtio_core_outputs_record0_rec_payload_channel != main_rtio_core_outputs_record2_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_rec_payload_fine_ts != main_rtio_core_outputs_record2_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record0_rec_payload_address != main_rtio_core_outputs_record2_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference4 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_121 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_122;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference5 <= 1'd0;
	if ((main_rtio_core_outputs_record1_rec_payload_channel != main_rtio_core_outputs_record3_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record1_rec_payload_fine_ts != main_rtio_core_outputs_record3_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record1_rec_payload_address != main_rtio_core_outputs_record3_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference5 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_122 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_123;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference6 <= 1'd0;
	if ((main_rtio_core_outputs_record4_rec_payload_channel != main_rtio_core_outputs_record6_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_rec_payload_fine_ts != main_rtio_core_outputs_record6_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record4_rec_payload_address != main_rtio_core_outputs_record6_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference6 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_123 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_124;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference7 <= 1'd0;
	if ((main_rtio_core_outputs_record5_rec_payload_channel != main_rtio_core_outputs_record7_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record5_rec_payload_fine_ts != main_rtio_core_outputs_record7_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record5_rec_payload_address != main_rtio_core_outputs_record7_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference7 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_124 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_125;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference8 <= 1'd0;
	if ((main_rtio_core_outputs_record9_rec_payload_channel != main_rtio_core_outputs_record10_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record9_rec_payload_fine_ts != main_rtio_core_outputs_record10_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record9_rec_payload_address != main_rtio_core_outputs_record10_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference8 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_125 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_126;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference9 <= 1'd0;
	if ((main_rtio_core_outputs_record13_rec_payload_channel != main_rtio_core_outputs_record14_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record13_rec_payload_fine_ts != main_rtio_core_outputs_record14_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record13_rec_payload_address != main_rtio_core_outputs_record14_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference9 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_126 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_127;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference10 <= 1'd0;
	if ((main_rtio_core_outputs_record16_rec_payload_channel != main_rtio_core_outputs_record20_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record16_rec_payload_fine_ts != main_rtio_core_outputs_record20_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record16_rec_payload_address != main_rtio_core_outputs_record20_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference10 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_127 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_128;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference11 <= 1'd0;
	if ((main_rtio_core_outputs_record17_rec_payload_channel != main_rtio_core_outputs_record21_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record17_rec_payload_fine_ts != main_rtio_core_outputs_record21_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record17_rec_payload_address != main_rtio_core_outputs_record21_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference11 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_128 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_129;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference12 <= 1'd0;
	if ((main_rtio_core_outputs_record18_rec_payload_channel != main_rtio_core_outputs_record22_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record18_rec_payload_fine_ts != main_rtio_core_outputs_record22_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record18_rec_payload_address != main_rtio_core_outputs_record22_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference12 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_129 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_130;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference13 <= 1'd0;
	if ((main_rtio_core_outputs_record19_rec_payload_channel != main_rtio_core_outputs_record23_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record19_rec_payload_fine_ts != main_rtio_core_outputs_record23_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record19_rec_payload_address != main_rtio_core_outputs_record23_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference13 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_130 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_131;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference14 <= 1'd0;
	if ((main_rtio_core_outputs_record26_rec_payload_channel != main_rtio_core_outputs_record28_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record26_rec_payload_fine_ts != main_rtio_core_outputs_record28_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record26_rec_payload_address != main_rtio_core_outputs_record28_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference14 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_131 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_132;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference15 <= 1'd0;
	if ((main_rtio_core_outputs_record27_rec_payload_channel != main_rtio_core_outputs_record29_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record27_rec_payload_fine_ts != main_rtio_core_outputs_record29_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record27_rec_payload_address != main_rtio_core_outputs_record29_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference15 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_132 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_133;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference16 <= 1'd0;
	if ((main_rtio_core_outputs_record33_rec_payload_channel != main_rtio_core_outputs_record34_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record33_rec_payload_fine_ts != main_rtio_core_outputs_record34_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record33_rec_payload_address != main_rtio_core_outputs_record34_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference16 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_133 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_134;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference17 <= 1'd0;
	if ((main_rtio_core_outputs_record35_rec_payload_channel != main_rtio_core_outputs_record36_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record35_rec_payload_fine_ts != main_rtio_core_outputs_record36_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record35_rec_payload_address != main_rtio_core_outputs_record36_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference17 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_134 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_135;
// synthesis translate_on
always @(*) begin
	main_rtio_core_outputs_nondata_difference18 <= 1'd0;
	if ((main_rtio_core_outputs_record37_rec_payload_channel != main_rtio_core_outputs_record38_rec_payload_channel)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record37_rec_payload_fine_ts != main_rtio_core_outputs_record38_rec_payload_fine_ts)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
	if ((main_rtio_core_outputs_record37_rec_payload_address != main_rtio_core_outputs_record38_rec_payload_address)) begin
		main_rtio_core_outputs_nondata_difference18 <= 1'd1;
	end
// synthesis translate_off
	dummy_d_135 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_din = {main_rtio_core_inputs_record0_fifo_in_timestamp, main_rtio_core_inputs_record0_fifo_in_data};
assign {main_rtio_core_inputs_record0_fifo_out_timestamp, main_rtio_core_inputs_record0_fifo_out_data} = main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout;
assign main_rtio_core_inputs_record0_fifo_in_data = main_inout_8x0_inout_8x0_iinterface0_data;
assign main_rtio_core_inputs_record0_fifo_in_timestamp = {main_coarse_ts, main_inout_8x0_inout_8x0_iinterface0_fine_ts};
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_we = main_inout_8x0_inout_8x0_iinterface0_stb;
assign main_rtio_core_inputs_overflow_io0 = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_we & (~main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable));
assign main_rtio_core_inputs_blindtransfer0_i = main_rtio_core_inputs_overflow_io0;
assign main_rtio_core_inputs_selected0 = (main_rtio_core_cri_chan_sel[15:0] == 2'd3);
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_re = ((main_rtio_core_inputs_selected0 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow0));
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_din = {main_rtio_core_inputs_record1_fifo_in_timestamp, main_rtio_core_inputs_record1_fifo_in_data};
assign {main_rtio_core_inputs_record1_fifo_out_timestamp, main_rtio_core_inputs_record1_fifo_out_data} = main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout;
assign main_rtio_core_inputs_record1_fifo_in_data = main_inout_8x1_inout_8x1_iinterface1_data;
assign main_rtio_core_inputs_record1_fifo_in_timestamp = {main_coarse_ts, main_inout_8x1_inout_8x1_iinterface1_fine_ts};
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_we = main_inout_8x1_inout_8x1_iinterface1_stb;
assign main_rtio_core_inputs_overflow_io1 = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_we & (~main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable));
assign main_rtio_core_inputs_blindtransfer1_i = main_rtio_core_inputs_overflow_io1;
assign main_rtio_core_inputs_selected1 = (main_rtio_core_cri_chan_sel[15:0] == 3'd7);
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_re = ((main_rtio_core_inputs_selected1 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow1));
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_din = {main_rtio_core_inputs_record2_fifo_in_timestamp, main_rtio_core_inputs_record2_fifo_in_data};
assign {main_rtio_core_inputs_record2_fifo_out_timestamp, main_rtio_core_inputs_record2_fifo_out_data} = main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout;
assign main_rtio_core_inputs_record2_fifo_in_data = main_inout_8x2_inout_8x2_iinterface2_data;
assign main_rtio_core_inputs_record2_fifo_in_timestamp = {main_coarse_ts, main_inout_8x2_inout_8x2_iinterface2_fine_ts};
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_we = main_inout_8x2_inout_8x2_iinterface2_stb;
assign main_rtio_core_inputs_overflow_io2 = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_we & (~main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable));
assign main_rtio_core_inputs_blindtransfer2_i = main_rtio_core_inputs_overflow_io2;
assign main_rtio_core_inputs_selected2 = (main_rtio_core_cri_chan_sel[15:0] == 4'd11);
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_re = ((main_rtio_core_inputs_selected2 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow2));
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_din = {main_rtio_core_inputs_record3_fifo_in_timestamp, main_rtio_core_inputs_record3_fifo_in_data};
assign {main_rtio_core_inputs_record3_fifo_out_timestamp, main_rtio_core_inputs_record3_fifo_out_data} = main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout;
assign main_rtio_core_inputs_record3_fifo_in_data = main_inout_8x3_inout_8x3_iinterface3_data;
assign main_rtio_core_inputs_record3_fifo_in_timestamp = {main_coarse_ts, main_inout_8x3_inout_8x3_iinterface3_fine_ts};
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_we = main_inout_8x3_inout_8x3_iinterface3_stb;
assign main_rtio_core_inputs_overflow_io3 = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_we & (~main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable));
assign main_rtio_core_inputs_blindtransfer3_i = main_rtio_core_inputs_overflow_io3;
assign main_rtio_core_inputs_selected3 = (main_rtio_core_cri_chan_sel[15:0] == 4'd15);
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_re = ((main_rtio_core_inputs_selected3 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow3));
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_din = {main_rtio_core_inputs_record4_fifo_in_timestamp, main_rtio_core_inputs_record4_fifo_in_data};
assign {main_rtio_core_inputs_record4_fifo_out_timestamp, main_rtio_core_inputs_record4_fifo_out_data} = main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout;
assign main_rtio_core_inputs_record4_fifo_in_data = main_inout_8x4_inout_8x4_iinterface4_data;
assign main_rtio_core_inputs_record4_fifo_in_timestamp = {main_coarse_ts, main_inout_8x4_inout_8x4_iinterface4_fine_ts};
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_we = main_inout_8x4_inout_8x4_iinterface4_stb;
assign main_rtio_core_inputs_overflow_io4 = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_we & (~main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable));
assign main_rtio_core_inputs_blindtransfer4_i = main_rtio_core_inputs_overflow_io4;
assign main_rtio_core_inputs_selected4 = (main_rtio_core_cri_chan_sel[15:0] == 5'd16);
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_re = ((main_rtio_core_inputs_selected4 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow4));
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_din = {main_rtio_core_inputs_record5_fifo_in_timestamp, main_rtio_core_inputs_record5_fifo_in_data};
assign {main_rtio_core_inputs_record5_fifo_out_timestamp, main_rtio_core_inputs_record5_fifo_out_data} = main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout;
assign main_rtio_core_inputs_record5_fifo_in_data = main_inout_8x5_inout_8x5_iinterface5_data;
assign main_rtio_core_inputs_record5_fifo_in_timestamp = {main_coarse_ts, main_inout_8x5_inout_8x5_iinterface5_fine_ts};
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_we = main_inout_8x5_inout_8x5_iinterface5_stb;
assign main_rtio_core_inputs_overflow_io5 = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_we & (~main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable));
assign main_rtio_core_inputs_blindtransfer5_i = main_rtio_core_inputs_overflow_io5;
assign main_rtio_core_inputs_selected5 = (main_rtio_core_cri_chan_sel[15:0] == 5'd17);
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_re = ((main_rtio_core_inputs_selected5 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow5));
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_din = {main_rtio_core_inputs_record6_fifo_in_timestamp, main_rtio_core_inputs_record6_fifo_in_data};
assign {main_rtio_core_inputs_record6_fifo_out_timestamp, main_rtio_core_inputs_record6_fifo_out_data} = main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout;
assign main_rtio_core_inputs_record6_fifo_in_data = main_inout_8x6_inout_8x6_iinterface6_data;
assign main_rtio_core_inputs_record6_fifo_in_timestamp = {main_coarse_ts, main_inout_8x6_inout_8x6_iinterface6_fine_ts};
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_we = main_inout_8x6_inout_8x6_iinterface6_stb;
assign main_rtio_core_inputs_overflow_io6 = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_we & (~main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable));
assign main_rtio_core_inputs_blindtransfer6_i = main_rtio_core_inputs_overflow_io6;
assign main_rtio_core_inputs_selected6 = (main_rtio_core_cri_chan_sel[15:0] == 5'd18);
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_re = ((main_rtio_core_inputs_selected6 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow6));
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_din = {main_rtio_core_inputs_record7_fifo_in_data};
assign {main_rtio_core_inputs_record7_fifo_out_data} = main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout;
assign main_rtio_core_inputs_record7_fifo_in_data = main_spimaster0_iinterface0_data;
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_we = main_spimaster0_iinterface0_stb;
assign main_rtio_core_inputs_overflow_io7 = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_we & (~main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable));
assign main_rtio_core_inputs_blindtransfer7_i = main_rtio_core_inputs_overflow_io7;
assign main_rtio_core_inputs_selected7 = (main_rtio_core_cri_chan_sel[15:0] == 5'd22);
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_re = ((main_rtio_core_inputs_selected7 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow7));
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_din = {main_rtio_core_inputs_record8_fifo_in_data};
assign {main_rtio_core_inputs_record8_fifo_out_data} = main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout;
assign main_rtio_core_inputs_record8_fifo_in_data = main_spimaster1_iinterface1_data;
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_we = main_spimaster1_iinterface1_stb;
assign main_rtio_core_inputs_overflow_io8 = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_we & (~main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable));
assign main_rtio_core_inputs_blindtransfer8_i = main_rtio_core_inputs_overflow_io8;
assign main_rtio_core_inputs_selected8 = (main_rtio_core_cri_chan_sel[15:0] == 5'd23);
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_re = ((main_rtio_core_inputs_selected8 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow8));
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_din = {main_rtio_core_inputs_record9_fifo_in_data};
assign {main_rtio_core_inputs_record9_fifo_out_data} = main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout;
assign main_rtio_core_inputs_record9_fifo_in_data = main_spimaster2_iinterface2_data;
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_we = main_spimaster2_iinterface2_stb;
assign main_rtio_core_inputs_overflow_io9 = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_we & (~main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable));
assign main_rtio_core_inputs_blindtransfer9_i = main_rtio_core_inputs_overflow_io9;
assign main_rtio_core_inputs_selected9 = (main_rtio_core_cri_chan_sel[15:0] == 5'd24);
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_re = ((main_rtio_core_inputs_selected9 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow9));
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_din = {main_rtio_core_inputs_record10_fifo_in_data};
assign {main_rtio_core_inputs_record10_fifo_out_data} = main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout;
assign main_rtio_core_inputs_record10_fifo_in_data = main_spimaster3_iinterface3_data;
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_we = main_spimaster3_iinterface3_stb;
assign main_rtio_core_inputs_overflow_io10 = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_we & (~main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable));
assign main_rtio_core_inputs_blindtransfer10_i = main_rtio_core_inputs_overflow_io10;
assign main_rtio_core_inputs_selected10 = (main_rtio_core_cri_chan_sel[15:0] == 5'd25);
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_re = ((main_rtio_core_inputs_selected10 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow10));
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_din = {main_rtio_core_inputs_record11_fifo_in_data};
assign {main_rtio_core_inputs_record11_fifo_out_data} = main_rtio_core_inputs_asyncfifo11_asyncfifo11_dout;
assign main_rtio_core_inputs_record11_fifo_in_data = main_spimaster4_iinterface4_data;
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_we = main_spimaster4_iinterface4_stb;
assign main_rtio_core_inputs_overflow_io11 = (main_rtio_core_inputs_asyncfifo11_asyncfifo11_we & (~main_rtio_core_inputs_asyncfifo11_asyncfifo11_writable));
assign main_rtio_core_inputs_blindtransfer11_i = main_rtio_core_inputs_overflow_io11;
assign main_rtio_core_inputs_selected11 = (main_rtio_core_cri_chan_sel[15:0] == 5'd26);
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_re = ((main_rtio_core_inputs_selected11 & main_rtio_core_inputs_i_ack) & (~main_rtio_core_inputs_overflow11));
assign main_rtio_core_inputs_i_status_raw = builder_comb_rhs_array_muxed9;
assign main_rtio_core_inputs_asyncfifo0_graycounter0_ce = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable & main_rtio_core_inputs_asyncfifo0_asyncfifo0_we);
assign main_rtio_core_inputs_asyncfifo0_graycounter1_ce = (main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & main_rtio_core_inputs_asyncfifo0_asyncfifo0_re);
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_writable = (((main_rtio_core_inputs_asyncfifo0_graycounter0_q[9] == main_rtio_core_inputs_asyncfifo0_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo0_graycounter0_q[8] == main_rtio_core_inputs_asyncfifo0_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo0_graycounter0_q[7:0] != main_rtio_core_inputs_asyncfifo0_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable = (main_rtio_core_inputs_asyncfifo0_graycounter1_q != main_rtio_core_inputs_asyncfifo0_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo0_wrport_adr = main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo0_wrport_dat_w = main_rtio_core_inputs_asyncfifo0_asyncfifo0_din;
assign main_rtio_core_inputs_asyncfifo0_wrport_we = main_rtio_core_inputs_asyncfifo0_graycounter0_ce;
assign main_rtio_core_inputs_asyncfifo0_rdport_adr = main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo0_asyncfifo0_dout = main_rtio_core_inputs_asyncfifo0_rdport_dat_r;

// synthesis translate_off
reg dummy_d_136;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo0_graycounter0_ce) begin
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= (main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary;
	end
// synthesis translate_off
	dummy_d_136 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_graycounter0_q_next = (main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary ^ main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_137;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo0_graycounter1_ce) begin
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= (main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary;
	end
// synthesis translate_off
	dummy_d_137 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo0_graycounter1_q_next = (main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary ^ main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer0_ps_i = (main_rtio_core_inputs_blindtransfer0_i & (~main_rtio_core_inputs_blindtransfer0_blind));
assign main_rtio_core_inputs_blindtransfer0_ps_ack_i = main_rtio_core_inputs_blindtransfer0_ps_o;
assign main_rtio_core_inputs_blindtransfer0_o = main_rtio_core_inputs_blindtransfer0_ps_o;
assign main_rtio_core_inputs_blindtransfer0_ps_o = (main_rtio_core_inputs_blindtransfer0_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer0_ps_ack_o = (main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo1_graycounter2_ce = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable & main_rtio_core_inputs_asyncfifo1_asyncfifo1_we);
assign main_rtio_core_inputs_asyncfifo1_graycounter3_ce = (main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & main_rtio_core_inputs_asyncfifo1_asyncfifo1_re);
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_writable = (((main_rtio_core_inputs_asyncfifo1_graycounter2_q[9] == main_rtio_core_inputs_asyncfifo1_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo1_graycounter2_q[8] == main_rtio_core_inputs_asyncfifo1_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo1_graycounter2_q[7:0] != main_rtio_core_inputs_asyncfifo1_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable = (main_rtio_core_inputs_asyncfifo1_graycounter3_q != main_rtio_core_inputs_asyncfifo1_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo1_wrport_adr = main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo1_wrport_dat_w = main_rtio_core_inputs_asyncfifo1_asyncfifo1_din;
assign main_rtio_core_inputs_asyncfifo1_wrport_we = main_rtio_core_inputs_asyncfifo1_graycounter2_ce;
assign main_rtio_core_inputs_asyncfifo1_rdport_adr = main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo1_asyncfifo1_dout = main_rtio_core_inputs_asyncfifo1_rdport_dat_r;

// synthesis translate_off
reg dummy_d_138;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo1_graycounter2_ce) begin
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= (main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary;
	end
// synthesis translate_off
	dummy_d_138 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo1_graycounter2_q_next = (main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary ^ main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_139;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo1_graycounter3_ce) begin
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= (main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary;
	end
// synthesis translate_off
	dummy_d_139 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo1_graycounter3_q_next = (main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary ^ main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer1_ps_i = (main_rtio_core_inputs_blindtransfer1_i & (~main_rtio_core_inputs_blindtransfer1_blind));
assign main_rtio_core_inputs_blindtransfer1_ps_ack_i = main_rtio_core_inputs_blindtransfer1_ps_o;
assign main_rtio_core_inputs_blindtransfer1_o = main_rtio_core_inputs_blindtransfer1_ps_o;
assign main_rtio_core_inputs_blindtransfer1_ps_o = (main_rtio_core_inputs_blindtransfer1_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer1_ps_ack_o = (main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo2_graycounter4_ce = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable & main_rtio_core_inputs_asyncfifo2_asyncfifo2_we);
assign main_rtio_core_inputs_asyncfifo2_graycounter5_ce = (main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & main_rtio_core_inputs_asyncfifo2_asyncfifo2_re);
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_writable = (((main_rtio_core_inputs_asyncfifo2_graycounter4_q[9] == main_rtio_core_inputs_asyncfifo2_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo2_graycounter4_q[8] == main_rtio_core_inputs_asyncfifo2_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo2_graycounter4_q[7:0] != main_rtio_core_inputs_asyncfifo2_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable = (main_rtio_core_inputs_asyncfifo2_graycounter5_q != main_rtio_core_inputs_asyncfifo2_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo2_wrport_adr = main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo2_wrport_dat_w = main_rtio_core_inputs_asyncfifo2_asyncfifo2_din;
assign main_rtio_core_inputs_asyncfifo2_wrport_we = main_rtio_core_inputs_asyncfifo2_graycounter4_ce;
assign main_rtio_core_inputs_asyncfifo2_rdport_adr = main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo2_asyncfifo2_dout = main_rtio_core_inputs_asyncfifo2_rdport_dat_r;

// synthesis translate_off
reg dummy_d_140;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo2_graycounter4_ce) begin
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= (main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary;
	end
// synthesis translate_off
	dummy_d_140 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo2_graycounter4_q_next = (main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary ^ main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_141;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo2_graycounter5_ce) begin
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= (main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary;
	end
// synthesis translate_off
	dummy_d_141 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo2_graycounter5_q_next = (main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary ^ main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer2_ps_i = (main_rtio_core_inputs_blindtransfer2_i & (~main_rtio_core_inputs_blindtransfer2_blind));
assign main_rtio_core_inputs_blindtransfer2_ps_ack_i = main_rtio_core_inputs_blindtransfer2_ps_o;
assign main_rtio_core_inputs_blindtransfer2_o = main_rtio_core_inputs_blindtransfer2_ps_o;
assign main_rtio_core_inputs_blindtransfer2_ps_o = (main_rtio_core_inputs_blindtransfer2_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer2_ps_ack_o = (main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo3_graycounter6_ce = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable & main_rtio_core_inputs_asyncfifo3_asyncfifo3_we);
assign main_rtio_core_inputs_asyncfifo3_graycounter7_ce = (main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & main_rtio_core_inputs_asyncfifo3_asyncfifo3_re);
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_writable = (((main_rtio_core_inputs_asyncfifo3_graycounter6_q[9] == main_rtio_core_inputs_asyncfifo3_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo3_graycounter6_q[8] == main_rtio_core_inputs_asyncfifo3_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo3_graycounter6_q[7:0] != main_rtio_core_inputs_asyncfifo3_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable = (main_rtio_core_inputs_asyncfifo3_graycounter7_q != main_rtio_core_inputs_asyncfifo3_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo3_wrport_adr = main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo3_wrport_dat_w = main_rtio_core_inputs_asyncfifo3_asyncfifo3_din;
assign main_rtio_core_inputs_asyncfifo3_wrport_we = main_rtio_core_inputs_asyncfifo3_graycounter6_ce;
assign main_rtio_core_inputs_asyncfifo3_rdport_adr = main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo3_asyncfifo3_dout = main_rtio_core_inputs_asyncfifo3_rdport_dat_r;

// synthesis translate_off
reg dummy_d_142;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo3_graycounter6_ce) begin
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= (main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary;
	end
// synthesis translate_off
	dummy_d_142 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo3_graycounter6_q_next = (main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary ^ main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_143;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo3_graycounter7_ce) begin
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= (main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary;
	end
// synthesis translate_off
	dummy_d_143 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo3_graycounter7_q_next = (main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary ^ main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer3_ps_i = (main_rtio_core_inputs_blindtransfer3_i & (~main_rtio_core_inputs_blindtransfer3_blind));
assign main_rtio_core_inputs_blindtransfer3_ps_ack_i = main_rtio_core_inputs_blindtransfer3_ps_o;
assign main_rtio_core_inputs_blindtransfer3_o = main_rtio_core_inputs_blindtransfer3_ps_o;
assign main_rtio_core_inputs_blindtransfer3_ps_o = (main_rtio_core_inputs_blindtransfer3_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer3_ps_ack_o = (main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo4_graycounter8_ce = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable & main_rtio_core_inputs_asyncfifo4_asyncfifo4_we);
assign main_rtio_core_inputs_asyncfifo4_graycounter9_ce = (main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & main_rtio_core_inputs_asyncfifo4_asyncfifo4_re);
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_writable = (((main_rtio_core_inputs_asyncfifo4_graycounter8_q[9] == main_rtio_core_inputs_asyncfifo4_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo4_graycounter8_q[8] == main_rtio_core_inputs_asyncfifo4_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo4_graycounter8_q[7:0] != main_rtio_core_inputs_asyncfifo4_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable = (main_rtio_core_inputs_asyncfifo4_graycounter9_q != main_rtio_core_inputs_asyncfifo4_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo4_wrport_adr = main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo4_wrport_dat_w = main_rtio_core_inputs_asyncfifo4_asyncfifo4_din;
assign main_rtio_core_inputs_asyncfifo4_wrport_we = main_rtio_core_inputs_asyncfifo4_graycounter8_ce;
assign main_rtio_core_inputs_asyncfifo4_rdport_adr = main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo4_asyncfifo4_dout = main_rtio_core_inputs_asyncfifo4_rdport_dat_r;

// synthesis translate_off
reg dummy_d_144;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo4_graycounter8_ce) begin
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= (main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary;
	end
// synthesis translate_off
	dummy_d_144 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo4_graycounter8_q_next = (main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary ^ main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_145;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo4_graycounter9_ce) begin
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= (main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary;
	end
// synthesis translate_off
	dummy_d_145 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo4_graycounter9_q_next = (main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary ^ main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer4_ps_i = (main_rtio_core_inputs_blindtransfer4_i & (~main_rtio_core_inputs_blindtransfer4_blind));
assign main_rtio_core_inputs_blindtransfer4_ps_ack_i = main_rtio_core_inputs_blindtransfer4_ps_o;
assign main_rtio_core_inputs_blindtransfer4_o = main_rtio_core_inputs_blindtransfer4_ps_o;
assign main_rtio_core_inputs_blindtransfer4_ps_o = (main_rtio_core_inputs_blindtransfer4_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer4_ps_ack_o = (main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo5_graycounter10_ce = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable & main_rtio_core_inputs_asyncfifo5_asyncfifo5_we);
assign main_rtio_core_inputs_asyncfifo5_graycounter11_ce = (main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & main_rtio_core_inputs_asyncfifo5_asyncfifo5_re);
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_writable = (((main_rtio_core_inputs_asyncfifo5_graycounter10_q[9] == main_rtio_core_inputs_asyncfifo5_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo5_graycounter10_q[8] == main_rtio_core_inputs_asyncfifo5_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo5_graycounter10_q[7:0] != main_rtio_core_inputs_asyncfifo5_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable = (main_rtio_core_inputs_asyncfifo5_graycounter11_q != main_rtio_core_inputs_asyncfifo5_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo5_wrport_adr = main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo5_wrport_dat_w = main_rtio_core_inputs_asyncfifo5_asyncfifo5_din;
assign main_rtio_core_inputs_asyncfifo5_wrport_we = main_rtio_core_inputs_asyncfifo5_graycounter10_ce;
assign main_rtio_core_inputs_asyncfifo5_rdport_adr = main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo5_asyncfifo5_dout = main_rtio_core_inputs_asyncfifo5_rdport_dat_r;

// synthesis translate_off
reg dummy_d_146;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo5_graycounter10_ce) begin
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= (main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary;
	end
// synthesis translate_off
	dummy_d_146 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo5_graycounter10_q_next = (main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary ^ main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_147;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo5_graycounter11_ce) begin
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= (main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary;
	end
// synthesis translate_off
	dummy_d_147 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo5_graycounter11_q_next = (main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary ^ main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer5_ps_i = (main_rtio_core_inputs_blindtransfer5_i & (~main_rtio_core_inputs_blindtransfer5_blind));
assign main_rtio_core_inputs_blindtransfer5_ps_ack_i = main_rtio_core_inputs_blindtransfer5_ps_o;
assign main_rtio_core_inputs_blindtransfer5_o = main_rtio_core_inputs_blindtransfer5_ps_o;
assign main_rtio_core_inputs_blindtransfer5_ps_o = (main_rtio_core_inputs_blindtransfer5_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer5_ps_ack_o = (main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo6_graycounter12_ce = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable & main_rtio_core_inputs_asyncfifo6_asyncfifo6_we);
assign main_rtio_core_inputs_asyncfifo6_graycounter13_ce = (main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & main_rtio_core_inputs_asyncfifo6_asyncfifo6_re);
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_writable = (((main_rtio_core_inputs_asyncfifo6_graycounter12_q[9] == main_rtio_core_inputs_asyncfifo6_consume_wdomain[9]) | (main_rtio_core_inputs_asyncfifo6_graycounter12_q[8] == main_rtio_core_inputs_asyncfifo6_consume_wdomain[8])) | (main_rtio_core_inputs_asyncfifo6_graycounter12_q[7:0] != main_rtio_core_inputs_asyncfifo6_consume_wdomain[7:0]));
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable = (main_rtio_core_inputs_asyncfifo6_graycounter13_q != main_rtio_core_inputs_asyncfifo6_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo6_wrport_adr = main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary[8:0];
assign main_rtio_core_inputs_asyncfifo6_wrport_dat_w = main_rtio_core_inputs_asyncfifo6_asyncfifo6_din;
assign main_rtio_core_inputs_asyncfifo6_wrport_we = main_rtio_core_inputs_asyncfifo6_graycounter12_ce;
assign main_rtio_core_inputs_asyncfifo6_rdport_adr = main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[8:0];
assign main_rtio_core_inputs_asyncfifo6_asyncfifo6_dout = main_rtio_core_inputs_asyncfifo6_rdport_dat_r;

// synthesis translate_off
reg dummy_d_148;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo6_graycounter12_ce) begin
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= (main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary;
	end
// synthesis translate_off
	dummy_d_148 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo6_graycounter12_q_next = (main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary ^ main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary[9:1]);

// synthesis translate_off
reg dummy_d_149;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= 10'd0;
	if (main_rtio_core_inputs_asyncfifo6_graycounter13_ce) begin
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= (main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary;
	end
// synthesis translate_off
	dummy_d_149 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo6_graycounter13_q_next = (main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary ^ main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary[9:1]);
assign main_rtio_core_inputs_blindtransfer6_ps_i = (main_rtio_core_inputs_blindtransfer6_i & (~main_rtio_core_inputs_blindtransfer6_blind));
assign main_rtio_core_inputs_blindtransfer6_ps_ack_i = main_rtio_core_inputs_blindtransfer6_ps_o;
assign main_rtio_core_inputs_blindtransfer6_o = main_rtio_core_inputs_blindtransfer6_ps_o;
assign main_rtio_core_inputs_blindtransfer6_ps_o = (main_rtio_core_inputs_blindtransfer6_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer6_ps_ack_o = (main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo7_graycounter14_ce = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable & main_rtio_core_inputs_asyncfifo7_asyncfifo7_we);
assign main_rtio_core_inputs_asyncfifo7_graycounter15_ce = (main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable & main_rtio_core_inputs_asyncfifo7_asyncfifo7_re);
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_writable = (((main_rtio_core_inputs_asyncfifo7_graycounter14_q[2] == main_rtio_core_inputs_asyncfifo7_consume_wdomain[2]) | (main_rtio_core_inputs_asyncfifo7_graycounter14_q[1] == main_rtio_core_inputs_asyncfifo7_consume_wdomain[1])) | (main_rtio_core_inputs_asyncfifo7_graycounter14_q[0] != main_rtio_core_inputs_asyncfifo7_consume_wdomain[0]));
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable = (main_rtio_core_inputs_asyncfifo7_graycounter15_q != main_rtio_core_inputs_asyncfifo7_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo7_wrport_adr = main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary[1:0];
assign main_rtio_core_inputs_asyncfifo7_wrport_dat_w = main_rtio_core_inputs_asyncfifo7_asyncfifo7_din;
assign main_rtio_core_inputs_asyncfifo7_wrport_we = main_rtio_core_inputs_asyncfifo7_graycounter14_ce;
assign main_rtio_core_inputs_asyncfifo7_rdport_adr = main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary[1:0];
assign main_rtio_core_inputs_asyncfifo7_asyncfifo7_dout = main_rtio_core_inputs_asyncfifo7_rdport_dat_r;

// synthesis translate_off
reg dummy_d_150;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo7_graycounter14_ce) begin
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= (main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary;
	end
// synthesis translate_off
	dummy_d_150 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo7_graycounter14_q_next = (main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary ^ main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_151;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo7_graycounter15_ce) begin
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= (main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary;
	end
// synthesis translate_off
	dummy_d_151 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo7_graycounter15_q_next = (main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary ^ main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary[2:1]);
assign main_rtio_core_inputs_blindtransfer7_ps_i = (main_rtio_core_inputs_blindtransfer7_i & (~main_rtio_core_inputs_blindtransfer7_blind));
assign main_rtio_core_inputs_blindtransfer7_ps_ack_i = main_rtio_core_inputs_blindtransfer7_ps_o;
assign main_rtio_core_inputs_blindtransfer7_o = main_rtio_core_inputs_blindtransfer7_ps_o;
assign main_rtio_core_inputs_blindtransfer7_ps_o = (main_rtio_core_inputs_blindtransfer7_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer7_ps_ack_o = (main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo8_graycounter16_ce = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable & main_rtio_core_inputs_asyncfifo8_asyncfifo8_we);
assign main_rtio_core_inputs_asyncfifo8_graycounter17_ce = (main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable & main_rtio_core_inputs_asyncfifo8_asyncfifo8_re);
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_writable = (((main_rtio_core_inputs_asyncfifo8_graycounter16_q[7] == main_rtio_core_inputs_asyncfifo8_consume_wdomain[7]) | (main_rtio_core_inputs_asyncfifo8_graycounter16_q[6] == main_rtio_core_inputs_asyncfifo8_consume_wdomain[6])) | (main_rtio_core_inputs_asyncfifo8_graycounter16_q[5:0] != main_rtio_core_inputs_asyncfifo8_consume_wdomain[5:0]));
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable = (main_rtio_core_inputs_asyncfifo8_graycounter17_q != main_rtio_core_inputs_asyncfifo8_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo8_wrport_adr = main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary[6:0];
assign main_rtio_core_inputs_asyncfifo8_wrport_dat_w = main_rtio_core_inputs_asyncfifo8_asyncfifo8_din;
assign main_rtio_core_inputs_asyncfifo8_wrport_we = main_rtio_core_inputs_asyncfifo8_graycounter16_ce;
assign main_rtio_core_inputs_asyncfifo8_rdport_adr = main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary[6:0];
assign main_rtio_core_inputs_asyncfifo8_asyncfifo8_dout = main_rtio_core_inputs_asyncfifo8_rdport_dat_r;

// synthesis translate_off
reg dummy_d_152;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo8_graycounter16_ce) begin
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= (main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary;
	end
// synthesis translate_off
	dummy_d_152 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo8_graycounter16_q_next = (main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary ^ main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_153;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo8_graycounter17_ce) begin
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= (main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary;
	end
// synthesis translate_off
	dummy_d_153 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo8_graycounter17_q_next = (main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary ^ main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary[7:1]);
assign main_rtio_core_inputs_blindtransfer8_ps_i = (main_rtio_core_inputs_blindtransfer8_i & (~main_rtio_core_inputs_blindtransfer8_blind));
assign main_rtio_core_inputs_blindtransfer8_ps_ack_i = main_rtio_core_inputs_blindtransfer8_ps_o;
assign main_rtio_core_inputs_blindtransfer8_o = main_rtio_core_inputs_blindtransfer8_ps_o;
assign main_rtio_core_inputs_blindtransfer8_ps_o = (main_rtio_core_inputs_blindtransfer8_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer8_ps_ack_o = (main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo9_graycounter18_ce = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable & main_rtio_core_inputs_asyncfifo9_asyncfifo9_we);
assign main_rtio_core_inputs_asyncfifo9_graycounter19_ce = (main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable & main_rtio_core_inputs_asyncfifo9_asyncfifo9_re);
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_writable = (((main_rtio_core_inputs_asyncfifo9_graycounter18_q[7] == main_rtio_core_inputs_asyncfifo9_consume_wdomain[7]) | (main_rtio_core_inputs_asyncfifo9_graycounter18_q[6] == main_rtio_core_inputs_asyncfifo9_consume_wdomain[6])) | (main_rtio_core_inputs_asyncfifo9_graycounter18_q[5:0] != main_rtio_core_inputs_asyncfifo9_consume_wdomain[5:0]));
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable = (main_rtio_core_inputs_asyncfifo9_graycounter19_q != main_rtio_core_inputs_asyncfifo9_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo9_wrport_adr = main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary[6:0];
assign main_rtio_core_inputs_asyncfifo9_wrport_dat_w = main_rtio_core_inputs_asyncfifo9_asyncfifo9_din;
assign main_rtio_core_inputs_asyncfifo9_wrport_we = main_rtio_core_inputs_asyncfifo9_graycounter18_ce;
assign main_rtio_core_inputs_asyncfifo9_rdport_adr = main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary[6:0];
assign main_rtio_core_inputs_asyncfifo9_asyncfifo9_dout = main_rtio_core_inputs_asyncfifo9_rdport_dat_r;

// synthesis translate_off
reg dummy_d_154;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo9_graycounter18_ce) begin
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= (main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary;
	end
// synthesis translate_off
	dummy_d_154 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo9_graycounter18_q_next = (main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary ^ main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_155;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo9_graycounter19_ce) begin
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= (main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary;
	end
// synthesis translate_off
	dummy_d_155 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo9_graycounter19_q_next = (main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary ^ main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary[7:1]);
assign main_rtio_core_inputs_blindtransfer9_ps_i = (main_rtio_core_inputs_blindtransfer9_i & (~main_rtio_core_inputs_blindtransfer9_blind));
assign main_rtio_core_inputs_blindtransfer9_ps_ack_i = main_rtio_core_inputs_blindtransfer9_ps_o;
assign main_rtio_core_inputs_blindtransfer9_o = main_rtio_core_inputs_blindtransfer9_ps_o;
assign main_rtio_core_inputs_blindtransfer9_ps_o = (main_rtio_core_inputs_blindtransfer9_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer9_ps_ack_o = (main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo10_graycounter20_ce = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable & main_rtio_core_inputs_asyncfifo10_asyncfifo10_we);
assign main_rtio_core_inputs_asyncfifo10_graycounter21_ce = (main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable & main_rtio_core_inputs_asyncfifo10_asyncfifo10_re);
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_writable = (((main_rtio_core_inputs_asyncfifo10_graycounter20_q[7] == main_rtio_core_inputs_asyncfifo10_consume_wdomain[7]) | (main_rtio_core_inputs_asyncfifo10_graycounter20_q[6] == main_rtio_core_inputs_asyncfifo10_consume_wdomain[6])) | (main_rtio_core_inputs_asyncfifo10_graycounter20_q[5:0] != main_rtio_core_inputs_asyncfifo10_consume_wdomain[5:0]));
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable = (main_rtio_core_inputs_asyncfifo10_graycounter21_q != main_rtio_core_inputs_asyncfifo10_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo10_wrport_adr = main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary[6:0];
assign main_rtio_core_inputs_asyncfifo10_wrport_dat_w = main_rtio_core_inputs_asyncfifo10_asyncfifo10_din;
assign main_rtio_core_inputs_asyncfifo10_wrport_we = main_rtio_core_inputs_asyncfifo10_graycounter20_ce;
assign main_rtio_core_inputs_asyncfifo10_rdport_adr = main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary[6:0];
assign main_rtio_core_inputs_asyncfifo10_asyncfifo10_dout = main_rtio_core_inputs_asyncfifo10_rdport_dat_r;

// synthesis translate_off
reg dummy_d_156;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo10_graycounter20_ce) begin
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= (main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary;
	end
// synthesis translate_off
	dummy_d_156 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo10_graycounter20_q_next = (main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary ^ main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary[7:1]);

// synthesis translate_off
reg dummy_d_157;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= 8'd0;
	if (main_rtio_core_inputs_asyncfifo10_graycounter21_ce) begin
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= (main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary;
	end
// synthesis translate_off
	dummy_d_157 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo10_graycounter21_q_next = (main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary ^ main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary[7:1]);
assign main_rtio_core_inputs_blindtransfer10_ps_i = (main_rtio_core_inputs_blindtransfer10_i & (~main_rtio_core_inputs_blindtransfer10_blind));
assign main_rtio_core_inputs_blindtransfer10_ps_ack_i = main_rtio_core_inputs_blindtransfer10_ps_o;
assign main_rtio_core_inputs_blindtransfer10_o = main_rtio_core_inputs_blindtransfer10_ps_o;
assign main_rtio_core_inputs_blindtransfer10_ps_o = (main_rtio_core_inputs_blindtransfer10_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer10_ps_ack_o = (main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r);
assign main_rtio_core_inputs_asyncfifo11_graycounter22_ce = (main_rtio_core_inputs_asyncfifo11_asyncfifo11_writable & main_rtio_core_inputs_asyncfifo11_asyncfifo11_we);
assign main_rtio_core_inputs_asyncfifo11_graycounter23_ce = (main_rtio_core_inputs_asyncfifo11_asyncfifo11_readable & main_rtio_core_inputs_asyncfifo11_asyncfifo11_re);
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_writable = (((main_rtio_core_inputs_asyncfifo11_graycounter22_q[2] == main_rtio_core_inputs_asyncfifo11_consume_wdomain[2]) | (main_rtio_core_inputs_asyncfifo11_graycounter22_q[1] == main_rtio_core_inputs_asyncfifo11_consume_wdomain[1])) | (main_rtio_core_inputs_asyncfifo11_graycounter22_q[0] != main_rtio_core_inputs_asyncfifo11_consume_wdomain[0]));
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_readable = (main_rtio_core_inputs_asyncfifo11_graycounter23_q != main_rtio_core_inputs_asyncfifo11_produce_rdomain);
assign main_rtio_core_inputs_asyncfifo11_wrport_adr = main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary[1:0];
assign main_rtio_core_inputs_asyncfifo11_wrport_dat_w = main_rtio_core_inputs_asyncfifo11_asyncfifo11_din;
assign main_rtio_core_inputs_asyncfifo11_wrport_we = main_rtio_core_inputs_asyncfifo11_graycounter22_ce;
assign main_rtio_core_inputs_asyncfifo11_rdport_adr = main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary[1:0];
assign main_rtio_core_inputs_asyncfifo11_asyncfifo11_dout = main_rtio_core_inputs_asyncfifo11_rdport_dat_r;

// synthesis translate_off
reg dummy_d_158;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo11_graycounter22_ce) begin
		main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary <= (main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary <= main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary;
	end
// synthesis translate_off
	dummy_d_158 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo11_graycounter22_q_next = (main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary ^ main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary[2:1]);

// synthesis translate_off
reg dummy_d_159;
// synthesis translate_on
always @(*) begin
	main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary <= 3'd0;
	if (main_rtio_core_inputs_asyncfifo11_graycounter23_ce) begin
		main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary <= (main_rtio_core_inputs_asyncfifo11_graycounter23_q_binary + 1'd1);
	end else begin
		main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary <= main_rtio_core_inputs_asyncfifo11_graycounter23_q_binary;
	end
// synthesis translate_off
	dummy_d_159 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_core_inputs_asyncfifo11_graycounter23_q_next = (main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary ^ main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary[2:1]);
assign main_rtio_core_inputs_blindtransfer11_ps_i = (main_rtio_core_inputs_blindtransfer11_i & (~main_rtio_core_inputs_blindtransfer11_blind));
assign main_rtio_core_inputs_blindtransfer11_ps_ack_i = main_rtio_core_inputs_blindtransfer11_ps_o;
assign main_rtio_core_inputs_blindtransfer11_o = main_rtio_core_inputs_blindtransfer11_ps_o;
assign main_rtio_core_inputs_blindtransfer11_ps_o = (main_rtio_core_inputs_blindtransfer11_ps_toggle_o ^ main_rtio_core_inputs_blindtransfer11_ps_toggle_o_r);
assign main_rtio_core_inputs_blindtransfer11_ps_ack_o = (main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o ^ main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o_r);
assign main_rtio_core_o_collision_sync_ps_i = (main_rtio_core_o_collision_sync_i & (~main_rtio_core_o_collision_sync_blind));
assign main_rtio_core_o_collision_sync_ps_ack_i = main_rtio_core_o_collision_sync_ps_o;
assign main_rtio_core_o_collision_sync_o = main_rtio_core_o_collision_sync_ps_o;
assign main_rtio_core_o_collision_sync_ps_o = (main_rtio_core_o_collision_sync_ps_toggle_o ^ main_rtio_core_o_collision_sync_ps_toggle_o_r);
assign main_rtio_core_o_collision_sync_ps_ack_o = (main_rtio_core_o_collision_sync_ps_ack_toggle_o ^ main_rtio_core_o_collision_sync_ps_ack_toggle_o_r);
assign main_rtio_core_o_busy_sync_ps_i = (main_rtio_core_o_busy_sync_i & (~main_rtio_core_o_busy_sync_blind));
assign main_rtio_core_o_busy_sync_ps_ack_i = main_rtio_core_o_busy_sync_ps_o;
assign main_rtio_core_o_busy_sync_o = main_rtio_core_o_busy_sync_ps_o;
assign main_rtio_core_o_busy_sync_ps_o = (main_rtio_core_o_busy_sync_ps_toggle_o ^ main_rtio_core_o_busy_sync_ps_toggle_o_r);
assign main_rtio_core_o_busy_sync_ps_ack_o = (main_rtio_core_o_busy_sync_ps_ack_toggle_o ^ main_rtio_core_o_busy_sync_ps_ack_toggle_o_r);
assign main_rtio_now_hi_w = main_rtio_now[63:32];
assign main_rtio_now_lo_w = main_rtio_now[31:0];

// synthesis translate_off
reg dummy_d_160;
// synthesis translate_on
always @(*) begin
	main_rtio_cri_cmd <= 2'd0;
	main_rtio_cri_cmd <= 1'd0;
	if (main_rtio_o_data_re) begin
		main_rtio_cri_cmd <= 1'd1;
	end
	if (main_rtio_i_timeout_re) begin
		main_rtio_cri_cmd <= 2'd2;
	end
// synthesis translate_off
	dummy_d_160 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_cri_chan_sel = main_rtio_target_storage[31:8];
assign main_rtio_cri_o_timestamp = main_rtio_now;
assign main_rtio_cri_o_data = main_rtio_o_data_storage;
assign main_rtio_cri_o_address = main_rtio_target_storage[7:0];
assign main_rtio_o_status_status = main_rtio_cri_o_status;
assign main_rtio_cri_i_timeout = main_rtio_i_timeout_storage;
assign main_rtio_i_data_status = main_rtio_cri_i_data;
assign main_rtio_i_timestamp_status = main_rtio_cri_i_timestamp;
assign main_rtio_i_status_status = main_rtio_cri_i_status;
assign main_rtio_o_data_dat_w = 1'd0;
assign main_rtio_o_data_we = main_rtio_target_re;
assign main_dma_rawslicer_sink_stb = main_dma_dma_source_stb;
assign main_dma_dma_source_ack = main_dma_rawslicer_sink_ack;
assign main_dma_rawslicer_sink_eop = main_dma_dma_source_eop;
assign main_dma_rawslicer_sink_payload_data = main_dma_dma_source_payload_data;
assign main_dma_time_offset_sink_stb = main_dma_record_converter_source_stb;
assign main_dma_record_converter_source_ack = main_dma_time_offset_sink_ack;
assign main_dma_time_offset_sink_eop = main_dma_record_converter_source_eop;
assign main_dma_time_offset_sink_payload_length = main_dma_record_converter_source_payload_length;
assign main_dma_time_offset_sink_payload_channel = main_dma_record_converter_source_payload_channel;
assign main_dma_time_offset_sink_payload_timestamp = main_dma_record_converter_source_payload_timestamp;
assign main_dma_time_offset_sink_payload_address = main_dma_record_converter_source_payload_address;
assign main_dma_time_offset_sink_payload_data = main_dma_record_converter_source_payload_data;
assign main_dma_cri_master_sink_stb = main_dma_time_offset_source_stb;
assign main_dma_time_offset_source_ack = main_dma_cri_master_sink_ack;
assign main_dma_cri_master_sink_eop = main_dma_time_offset_source_eop;
assign main_dma_cri_master_sink_payload_length = main_dma_time_offset_source_payload_length;
assign main_dma_cri_master_sink_payload_channel = main_dma_time_offset_source_payload_channel;
assign main_dma_cri_master_sink_payload_timestamp = main_dma_time_offset_source_payload_timestamp;
assign main_dma_cri_master_sink_payload_address = main_dma_time_offset_source_payload_address;
assign main_dma_cri_master_sink_payload_data = main_dma_time_offset_source_payload_data;
assign main_dma_dma_bus_stb = (main_dma_dma_sink_stb & ((~main_dma_dma_data_reg_loaded) | main_dma_dma_source_ack));
assign main_interface0_bus_cyc = main_dma_dma_bus_stb;
assign main_interface0_bus_stb = main_dma_dma_bus_stb;
assign main_interface0_bus_adr = main_dma_dma_sink_payload_address;
assign main_dma_dma_sink_ack = main_interface0_bus_ack;
assign main_dma_dma_source_stb = main_dma_dma_data_reg_loaded;
assign main_dma_rawslicer_source = main_dma_rawslicer_buf[615:0];

// synthesis translate_off
reg dummy_d_161;
// synthesis translate_on
always @(*) begin
	main_dma_rawslicer_sink_ack <= 1'd0;
	main_dma_rawslicer_source_stb <= 1'd0;
	main_dma_rawslicer_flush_done <= 1'd0;
	main_dma_rawslicer_next_level <= 8'd0;
	main_dma_rawslicer_load_buf <= 1'd0;
	main_dma_rawslicer_shift_buf <= 1'd0;
	builder_resetinserter_next_state <= 2'd0;
	main_dma_rawslicer_next_level <= main_dma_rawslicer_level;
	builder_resetinserter_next_state <= builder_resetinserter_state;
	case (builder_resetinserter_state)
		1'd1: begin
			main_dma_rawslicer_source_stb <= 1'd1;
			main_dma_rawslicer_shift_buf <= 1'd1;
			main_dma_rawslicer_next_level <= (main_dma_rawslicer_level - main_dma_rawslicer_source_consume);
			if ((main_dma_rawslicer_next_level < 7'd77)) begin
				builder_resetinserter_next_state <= 1'd0;
			end
			if (main_dma_rawslicer_flush) begin
				builder_resetinserter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_dma_rawslicer_next_level <= 1'd0;
			main_dma_rawslicer_sink_ack <= 1'd1;
			if ((main_dma_rawslicer_sink_stb & main_dma_rawslicer_sink_eop)) begin
				main_dma_rawslicer_flush_done <= 1'd1;
				builder_resetinserter_next_state <= 1'd0;
			end
		end
		default: begin
			main_dma_rawslicer_sink_ack <= 1'd1;
			main_dma_rawslicer_load_buf <= 1'd1;
			if (main_dma_rawslicer_sink_stb) begin
				main_dma_rawslicer_next_level <= (main_dma_rawslicer_level + 7'd64);
			end
			if ((main_dma_rawslicer_next_level >= 7'd77)) begin
				builder_resetinserter_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_161 <= dummy_s;
// synthesis translate_on
end
assign {main_dma_record_converter_record_raw_data, main_dma_record_converter_record_raw_address, main_dma_record_converter_record_raw_timestamp, main_dma_record_converter_record_raw_channel, main_dma_record_converter_record_raw_length} = main_dma_rawslicer_source;
assign main_dma_record_converter_source_payload_channel = main_dma_record_converter_record_raw_channel;
assign main_dma_record_converter_source_payload_timestamp = main_dma_record_converter_record_raw_timestamp;
assign main_dma_record_converter_source_payload_address = main_dma_record_converter_record_raw_address;

// synthesis translate_off
reg dummy_d_162;
// synthesis translate_on
always @(*) begin
	main_dma_record_converter_source_payload_data <= 512'd0;
	case (main_dma_record_converter_record_raw_length)
		4'd14: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[7:0];
		end
		4'd15: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[15:0];
		end
		5'd16: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[23:0];
		end
		5'd17: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[31:0];
		end
		5'd18: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[39:0];
		end
		5'd19: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[47:0];
		end
		5'd20: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[55:0];
		end
		5'd21: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[63:0];
		end
		5'd22: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[71:0];
		end
		5'd23: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[79:0];
		end
		5'd24: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[87:0];
		end
		5'd25: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[95:0];
		end
		5'd26: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[103:0];
		end
		5'd27: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[111:0];
		end
		5'd28: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[119:0];
		end
		5'd29: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[127:0];
		end
		5'd30: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[135:0];
		end
		5'd31: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[143:0];
		end
		6'd32: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[151:0];
		end
		6'd33: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[159:0];
		end
		6'd34: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[167:0];
		end
		6'd35: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[175:0];
		end
		6'd36: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[183:0];
		end
		6'd37: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[191:0];
		end
		6'd38: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[199:0];
		end
		6'd39: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[207:0];
		end
		6'd40: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[215:0];
		end
		6'd41: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[223:0];
		end
		6'd42: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[231:0];
		end
		6'd43: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[239:0];
		end
		6'd44: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[247:0];
		end
		6'd45: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[255:0];
		end
		6'd46: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[263:0];
		end
		6'd47: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[271:0];
		end
		6'd48: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[279:0];
		end
		6'd49: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[287:0];
		end
		6'd50: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[295:0];
		end
		6'd51: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[303:0];
		end
		6'd52: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[311:0];
		end
		6'd53: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[319:0];
		end
		6'd54: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[327:0];
		end
		6'd55: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[335:0];
		end
		6'd56: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[343:0];
		end
		6'd57: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[351:0];
		end
		6'd58: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[359:0];
		end
		6'd59: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[367:0];
		end
		6'd60: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[375:0];
		end
		6'd61: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[383:0];
		end
		6'd62: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[391:0];
		end
		6'd63: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[399:0];
		end
		7'd64: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[407:0];
		end
		7'd65: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[415:0];
		end
		7'd66: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[423:0];
		end
		7'd67: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[431:0];
		end
		7'd68: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[439:0];
		end
		7'd69: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[447:0];
		end
		7'd70: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[455:0];
		end
		7'd71: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[463:0];
		end
		7'd72: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[471:0];
		end
		7'd73: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[479:0];
		end
		7'd74: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[487:0];
		end
		7'd75: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[495:0];
		end
		7'd76: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[503:0];
		end
		7'd77: begin
			main_dma_record_converter_source_payload_data <= main_dma_record_converter_record_raw_data[511:0];
		end
	endcase
// synthesis translate_off
	dummy_d_162 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_163;
// synthesis translate_on
always @(*) begin
	main_dma_rawslicer_source_consume <= 7'd0;
	main_dma_rawslicer_flush <= 1'd0;
	main_dma_record_converter_source_stb <= 1'd0;
	main_dma_record_converter_source_eop <= 1'd0;
	main_dma_record_converter_end_marker_found <= 1'd0;
	builder_recordconverter_next_state <= 2'd0;
	builder_recordconverter_next_state <= builder_recordconverter_state;
	case (builder_recordconverter_state)
		1'd1: begin
			main_dma_record_converter_end_marker_found <= 1'd1;
			if (main_dma_record_converter_flush) begin
				main_dma_rawslicer_flush <= 1'd1;
				builder_recordconverter_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (main_dma_rawslicer_flush_done) begin
				builder_recordconverter_next_state <= 2'd3;
			end
		end
		2'd3: begin
			main_dma_record_converter_source_eop <= 1'd1;
			main_dma_record_converter_source_stb <= 1'd1;
			if (main_dma_record_converter_source_ack) begin
				builder_recordconverter_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_dma_rawslicer_source_stb) begin
				if ((main_dma_record_converter_record_raw_length == 1'd0)) begin
					builder_recordconverter_next_state <= 1'd1;
				end else begin
					main_dma_record_converter_source_stb <= 1'd1;
				end
			end
			if (main_dma_record_converter_source_ack) begin
				main_dma_rawslicer_source_consume <= main_dma_record_converter_record_raw_length;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_163 <= dummy_s;
// synthesis translate_on
end
assign main_dma_time_offset_sink_ack = (~main_dma_time_offset_source_stb);
assign main_dma_cri_master_cri_chan_sel = main_dma_cri_master_sink_payload_channel;
assign main_dma_cri_master_cri_o_timestamp = main_dma_cri_master_sink_payload_timestamp;
assign main_dma_cri_master_cri_o_address = main_dma_cri_master_sink_payload_address;
assign main_dma_cri_master_cri_o_data = main_dma_cri_master_sink_payload_data;

// synthesis translate_off
reg dummy_d_164;
// synthesis translate_on
always @(*) begin
	main_dma_cri_master_sink_ack <= 1'd0;
	main_dma_cri_master_cri_cmd <= 2'd0;
	main_dma_cri_master_busy <= 1'd0;
	main_dma_cri_master_underflow_trigger <= 1'd0;
	main_dma_cri_master_link_error_trigger <= 1'd0;
	builder_crimaster_next_state <= 3'd0;
	builder_crimaster_next_state <= builder_crimaster_state;
	case (builder_crimaster_state)
		1'd1: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_cri_cmd <= 1'd1;
			builder_crimaster_next_state <= 2'd2;
		end
		2'd2: begin
			main_dma_cri_master_busy <= 1'd1;
			if ((main_dma_cri_master_cri_o_status == 1'd0)) begin
				main_dma_cri_master_sink_ack <= 1'd1;
				builder_crimaster_next_state <= 1'd0;
			end
			if (main_dma_cri_master_cri_o_status[1]) begin
				builder_crimaster_next_state <= 2'd3;
			end
			if (main_dma_cri_master_cri_o_status[2]) begin
				builder_crimaster_next_state <= 3'd4;
			end
		end
		2'd3: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_underflow_trigger <= 1'd1;
			main_dma_cri_master_sink_ack <= 1'd1;
			builder_crimaster_next_state <= 1'd0;
		end
		3'd4: begin
			main_dma_cri_master_busy <= 1'd1;
			main_dma_cri_master_link_error_trigger <= 1'd1;
			main_dma_cri_master_sink_ack <= 1'd1;
			builder_crimaster_next_state <= 1'd0;
		end
		default: begin
			if ((main_dma_cri_master_error_w == 1'd0)) begin
				if (main_dma_cri_master_sink_stb) begin
					if (main_dma_cri_master_sink_eop) begin
						main_dma_cri_master_sink_ack <= 1'd1;
					end else begin
						builder_crimaster_next_state <= 1'd1;
					end
				end
			end else begin
				main_dma_cri_master_sink_ack <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_164 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_165;
// synthesis translate_on
always @(*) begin
	main_dma_enable_enable_w <= 1'd0;
	main_dma_flow_enable <= 1'd0;
	main_dma_record_converter_flush <= 1'd0;
	builder_fsm_next_state <= 3'd0;
	builder_fsm_next_state <= builder_fsm_state;
	case (builder_fsm_state)
		1'd1: begin
			main_dma_enable_enable_w <= 1'd1;
			main_dma_flow_enable <= 1'd1;
			if (main_dma_record_converter_end_marker_found) begin
				builder_fsm_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_dma_enable_enable_w <= 1'd1;
			main_dma_record_converter_flush <= 1'd1;
			builder_fsm_next_state <= 2'd3;
		end
		2'd3: begin
			main_dma_enable_enable_w <= 1'd1;
			if (((main_dma_cri_master_sink_stb & main_dma_cri_master_sink_ack) & main_dma_cri_master_sink_eop)) begin
				builder_fsm_next_state <= 3'd4;
			end
		end
		3'd4: begin
			main_dma_enable_enable_w <= 1'd1;
			if ((~main_dma_cri_master_busy)) begin
				builder_fsm_next_state <= 1'd0;
			end
		end
		default: begin
			if (main_dma_enable_enable_re) begin
				builder_fsm_next_state <= 1'd1;
			end
		end
	endcase
// synthesis translate_off
	dummy_d_165 <= dummy_s;
// synthesis translate_on
end
assign main_csrbank0_target0_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_target0_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 1'd0));
assign main_rtio_now_hi_r = main_csrbank0_bus_dat_w[31:0];
assign main_rtio_now_hi_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 1'd1));
assign main_rtio_now_lo_r = main_csrbank0_bus_dat_w[31:0];
assign main_rtio_now_lo_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 2'd2));
assign main_csrbank0_o_data15_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data15_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 2'd3));
assign main_csrbank0_o_data14_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data14_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 3'd4));
assign main_csrbank0_o_data13_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data13_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 3'd5));
assign main_csrbank0_o_data12_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data12_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 3'd6));
assign main_csrbank0_o_data11_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data11_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 3'd7));
assign main_csrbank0_o_data10_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data10_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd8));
assign main_csrbank0_o_data9_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data9_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd9));
assign main_csrbank0_o_data8_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data8_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd10));
assign main_csrbank0_o_data7_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data7_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd11));
assign main_csrbank0_o_data6_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data6_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd12));
assign main_csrbank0_o_data5_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data5_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd13));
assign main_csrbank0_o_data4_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data4_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd14));
assign main_csrbank0_o_data3_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data3_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 4'd15));
assign main_csrbank0_o_data2_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data2_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd16));
assign main_csrbank0_o_data1_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data1_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd17));
assign main_csrbank0_o_data0_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_o_data0_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd18));
assign main_csrbank0_o_status_r = main_csrbank0_bus_dat_w[2:0];
assign main_csrbank0_o_status_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd19));
assign main_csrbank0_i_timeout1_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_i_timeout1_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd20));
assign main_csrbank0_i_timeout0_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_i_timeout0_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd21));
assign main_csrbank0_i_data_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_i_data_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd22));
assign main_csrbank0_i_timestamp1_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_i_timestamp1_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd23));
assign main_csrbank0_i_timestamp0_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_i_timestamp0_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd24));
assign main_csrbank0_i_status_r = main_csrbank0_bus_dat_w[3:0];
assign main_csrbank0_i_status_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd25));
assign main_rtio_i_overflow_reset_r = main_csrbank0_bus_dat_w[0];
assign main_rtio_i_overflow_reset_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd26));
assign main_csrbank0_counter1_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_counter1_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd27));
assign main_csrbank0_counter0_r = main_csrbank0_bus_dat_w[31:0];
assign main_csrbank0_counter0_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd28));
assign main_rtio_counter_update_r = main_csrbank0_bus_dat_w[0];
assign main_rtio_counter_update_re = ((((main_csrbank0_bus_cyc & main_csrbank0_bus_stb) & (~main_csrbank0_bus_ack)) & main_csrbank0_bus_we) & (main_csrbank0_bus_adr[4:0] == 5'd29));
assign main_rtio_target_storage = main_rtio_target_storage_full[31:0];
assign main_csrbank0_target0_w = main_rtio_target_storage_full[31:0];
assign main_rtio_o_data_storage = main_rtio_o_data_storage_full[511:0];
assign main_csrbank0_o_data15_w = main_rtio_o_data_storage_full[511:480];
assign main_csrbank0_o_data14_w = main_rtio_o_data_storage_full[479:448];
assign main_csrbank0_o_data13_w = main_rtio_o_data_storage_full[447:416];
assign main_csrbank0_o_data12_w = main_rtio_o_data_storage_full[415:384];
assign main_csrbank0_o_data11_w = main_rtio_o_data_storage_full[383:352];
assign main_csrbank0_o_data10_w = main_rtio_o_data_storage_full[351:320];
assign main_csrbank0_o_data9_w = main_rtio_o_data_storage_full[319:288];
assign main_csrbank0_o_data8_w = main_rtio_o_data_storage_full[287:256];
assign main_csrbank0_o_data7_w = main_rtio_o_data_storage_full[255:224];
assign main_csrbank0_o_data6_w = main_rtio_o_data_storage_full[223:192];
assign main_csrbank0_o_data5_w = main_rtio_o_data_storage_full[191:160];
assign main_csrbank0_o_data4_w = main_rtio_o_data_storage_full[159:128];
assign main_csrbank0_o_data3_w = main_rtio_o_data_storage_full[127:96];
assign main_csrbank0_o_data2_w = main_rtio_o_data_storage_full[95:64];
assign main_csrbank0_o_data1_w = main_rtio_o_data_storage_full[63:32];
assign main_csrbank0_o_data0_w = main_rtio_o_data_storage_full[31:0];
assign main_csrbank0_o_status_w = main_rtio_o_status_status[2:0];
assign main_rtio_i_timeout_storage = main_rtio_i_timeout_storage_full[63:0];
assign main_csrbank0_i_timeout1_w = main_rtio_i_timeout_storage_full[63:32];
assign main_csrbank0_i_timeout0_w = main_rtio_i_timeout_storage_full[31:0];
assign main_csrbank0_i_data_w = main_rtio_i_data_status[31:0];
assign main_csrbank0_i_timestamp1_w = main_rtio_i_timestamp_status[63:32];
assign main_csrbank0_i_timestamp0_w = main_rtio_i_timestamp_status[31:0];
assign main_csrbank0_i_status_w = main_rtio_i_status_status[3:0];
assign main_csrbank0_counter1_w = main_rtio_counter_status[63:32];
assign main_csrbank0_counter0_w = main_rtio_counter_status[31:0];
assign main_dma_enable_enable_r = main_csrbank1_bus_dat_w[0];
assign main_dma_enable_enable_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 1'd0));
assign main_csrbank1_base_address1_r = main_csrbank1_bus_dat_w[3:0];
assign main_csrbank1_base_address1_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 1'd1));
assign main_csrbank1_base_address0_r = main_csrbank1_bus_dat_w[31:0];
assign main_csrbank1_base_address0_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 2'd2));
assign main_csrbank1_time_offset1_r = main_csrbank1_bus_dat_w[31:0];
assign main_csrbank1_time_offset1_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 2'd3));
assign main_csrbank1_time_offset0_r = main_csrbank1_bus_dat_w[31:0];
assign main_csrbank1_time_offset0_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 3'd4));
assign main_dma_cri_master_error_r = main_csrbank1_bus_dat_w[1:0];
assign main_dma_cri_master_error_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 3'd5));
assign main_csrbank1_error_channel_r = main_csrbank1_bus_dat_w[23:0];
assign main_csrbank1_error_channel_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 3'd6));
assign main_csrbank1_error_timestamp1_r = main_csrbank1_bus_dat_w[31:0];
assign main_csrbank1_error_timestamp1_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 3'd7));
assign main_csrbank1_error_timestamp0_r = main_csrbank1_bus_dat_w[31:0];
assign main_csrbank1_error_timestamp0_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 4'd8));
assign main_csrbank1_error_address_r = main_csrbank1_bus_dat_w[15:0];
assign main_csrbank1_error_address_re = ((((main_csrbank1_bus_cyc & main_csrbank1_bus_stb) & (~main_csrbank1_bus_ack)) & main_csrbank1_bus_we) & (main_csrbank1_bus_adr[3:0] == 4'd9));
assign main_dma_dma_storage = main_dma_dma_storage_full[35:6];
assign main_csrbank1_base_address1_w = main_dma_dma_storage_full[35:32];
assign main_csrbank1_base_address0_w = {main_dma_dma_storage_full[31:6], {26{1'd0}}};
assign main_dma_time_offset_storage = main_dma_time_offset_storage_full[63:0];
assign main_csrbank1_time_offset1_w = main_dma_time_offset_storage_full[63:32];
assign main_csrbank1_time_offset0_w = main_dma_time_offset_storage_full[31:0];
assign main_csrbank1_error_channel_w = main_dma_cri_master_error_channel_status[23:0];
assign main_csrbank1_error_timestamp1_w = main_dma_cri_master_error_timestamp_status[63:32];
assign main_csrbank1_error_timestamp0_w = main_dma_cri_master_error_timestamp_status[31:0];
assign main_csrbank1_error_address_w = main_dma_cri_master_error_address_status[15:0];
assign main_cri_con_shared_cmd = builder_comb_rhs_array_muxed10;
assign main_cri_con_shared_chan_sel = builder_comb_rhs_array_muxed11;
assign main_cri_con_shared_o_timestamp = builder_comb_rhs_array_muxed12;
assign main_cri_con_shared_o_data = builder_comb_rhs_array_muxed13;
assign main_cri_con_shared_o_address = builder_comb_rhs_array_muxed14;
assign main_cri_con_shared_i_timeout = builder_comb_rhs_array_muxed15;
assign main_rtio_cri_o_status = main_cri_con_shared_o_status;
assign main_dma_cri_master_cri_o_status = main_cri_con_shared_o_status;
assign main_rtio_cri_o_buffer_space_valid = main_cri_con_shared_o_buffer_space_valid;
assign main_dma_cri_master_cri_o_buffer_space_valid = main_cri_con_shared_o_buffer_space_valid;
assign main_rtio_cri_o_buffer_space = main_cri_con_shared_o_buffer_space;
assign main_dma_cri_master_cri_o_buffer_space = main_cri_con_shared_o_buffer_space;
assign main_rtio_cri_i_data = main_cri_con_shared_i_data;
assign main_dma_cri_master_cri_i_data = main_cri_con_shared_i_data;
assign main_rtio_cri_i_timestamp = main_cri_con_shared_i_timestamp;
assign main_dma_cri_master_cri_i_timestamp = main_cri_con_shared_i_timestamp;
assign main_rtio_cri_i_status = main_cri_con_shared_i_status;
assign main_dma_cri_master_cri_i_status = main_cri_con_shared_i_status;
assign main_rtio_core_cri_chan_sel = main_cri_con_shared_chan_sel;
assign main_rtio_core_cri_o_timestamp = main_cri_con_shared_o_timestamp;
assign main_rtio_core_cri_o_data = main_cri_con_shared_o_data;
assign main_rtio_core_cri_o_address = main_cri_con_shared_o_address;
assign main_rtio_core_cri_i_timeout = main_cri_con_shared_i_timeout;

// synthesis translate_off
reg dummy_d_166;
// synthesis translate_on
always @(*) begin
	main_rtio_core_cri_cmd <= 2'd0;
	if ((main_cri_con_selected == 1'd0)) begin
		main_rtio_core_cri_cmd <= main_cri_con_shared_cmd;
	end
// synthesis translate_off
	dummy_d_166 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_167;
// synthesis translate_on
always @(*) begin
	main_cri_con_shared_o_status <= 3'd0;
	main_cri_con_shared_o_buffer_space_valid <= 1'd0;
	main_cri_con_shared_o_buffer_space <= 16'd0;
	main_cri_con_shared_i_data <= 32'd0;
	main_cri_con_shared_i_timestamp <= 64'd0;
	main_cri_con_shared_i_status <= 4'd0;
	case (main_cri_con_selected)
		1'd0: begin
			main_cri_con_shared_o_status <= main_rtio_core_cri_o_status;
			main_cri_con_shared_o_buffer_space_valid <= main_rtio_core_cri_o_buffer_space_valid;
			main_cri_con_shared_o_buffer_space <= main_rtio_core_cri_o_buffer_space;
			main_cri_con_shared_i_data <= main_rtio_core_cri_i_data;
			main_cri_con_shared_i_timestamp <= main_rtio_core_cri_i_timestamp;
			main_cri_con_shared_i_status <= main_rtio_core_cri_i_status;
		end
	endcase
// synthesis translate_off
	dummy_d_167 <= dummy_s;
// synthesis translate_on
end
assign main_csrbank2_selected0_r = main_csrbank2_bus_dat_w[1:0];
assign main_csrbank2_selected0_re = ((((main_csrbank2_bus_cyc & main_csrbank2_bus_stb) & (~main_csrbank2_bus_ack)) & main_csrbank2_bus_we) & (main_csrbank2_bus_adr[0] == 1'd0));
assign main_cri_con_storage = main_cri_con_storage_full[1:0];
assign main_csrbank2_selected0_w = main_cri_con_storage_full[1:0];
assign main_mon_bussynchronizer0_i = main_output_8x0_o[7];
assign main_mon_bussynchronizer1_i = main_output_8x1_o[7];
assign main_mon_bussynchronizer2_i = main_output_8x2_o[7];
assign main_mon_bussynchronizer3_i = main_inout_8x0_serdes_i0[7];
assign main_mon_bussynchronizer4_i = main_inout_8x0_serdes_oe;
assign main_mon_bussynchronizer5_i = main_output_8x3_o[7];
assign main_mon_bussynchronizer6_i = main_output_8x4_o[7];
assign main_mon_bussynchronizer7_i = main_output_8x5_o[7];
assign main_mon_bussynchronizer8_i = main_inout_8x1_serdes_i0[7];
assign main_mon_bussynchronizer9_i = main_inout_8x1_serdes_oe;
assign main_mon_bussynchronizer10_i = main_output_8x6_o[7];
assign main_mon_bussynchronizer11_i = main_output_8x7_o[7];
assign main_mon_bussynchronizer12_i = main_output_8x8_o[7];
assign main_mon_bussynchronizer13_i = main_inout_8x2_serdes_i0[7];
assign main_mon_bussynchronizer14_i = main_inout_8x2_serdes_oe;
assign main_mon_bussynchronizer15_i = main_output_8x9_o[7];
assign main_mon_bussynchronizer16_i = main_output_8x10_o[7];
assign main_mon_bussynchronizer17_i = main_output_8x11_o[7];
assign main_mon_bussynchronizer18_i = main_inout_8x3_serdes_i0[7];
assign main_mon_bussynchronizer19_i = main_inout_8x3_serdes_oe;
assign main_mon_bussynchronizer20_i = main_inout_8x4_serdes_i0[7];
assign main_mon_bussynchronizer21_i = main_inout_8x4_serdes_oe;
assign main_mon_bussynchronizer22_i = main_inout_8x5_serdes_i0[7];
assign main_mon_bussynchronizer23_i = main_inout_8x5_serdes_oe;
assign main_mon_bussynchronizer24_i = main_inout_8x6_serdes_i0[7];
assign main_mon_bussynchronizer25_i = main_inout_8x6_serdes_oe;
assign main_mon_bussynchronizer26_i = main_output0_pad_o;
assign main_mon_bussynchronizer27_i = main_output1_pad_o;
assign main_mon_bussynchronizer28_i = main_ad9914_probes0;
assign main_mon_bussynchronizer29_i = main_ad9914_probes1;
assign main_mon_bussynchronizer30_i = main_ad9914_probes2;
assign main_mon_bussynchronizer31_i = main_ad9914_probes3;
assign main_mon_bussynchronizer32_i = main_ad9914_probes4;
assign main_mon_bussynchronizer33_i = main_ad9914_probes5;
assign main_mon_bussynchronizer34_i = main_ad9914_probes6;
assign main_mon_bussynchronizer35_i = main_ad9914_probes7;
assign main_mon_bussynchronizer36_i = main_ad9914_probes8;
assign main_mon_bussynchronizer37_i = main_ad9914_probes9;
assign main_mon_bussynchronizer38_i = main_ad9914_probes10;
assign main_mon_bussynchronizer28_wait = (~main_mon_bussynchronizer28_ping_i);
assign main_mon_bussynchronizer28_ping_i = ((main_mon_bussynchronizer28_starter | main_mon_bussynchronizer28_pong_o) | main_mon_bussynchronizer28_done);
assign main_mon_bussynchronizer28_pong_i = main_mon_bussynchronizer28_ping_o1;
assign main_mon_bussynchronizer28_ping_o0 = (main_mon_bussynchronizer28_ping_toggle_o ^ main_mon_bussynchronizer28_ping_toggle_o_r);
assign main_mon_bussynchronizer28_pong_o = (main_mon_bussynchronizer28_pong_toggle_o ^ main_mon_bussynchronizer28_pong_toggle_o_r);
assign main_mon_bussynchronizer28_done = (main_mon_bussynchronizer28_count == 1'd0);
assign main_mon_bussynchronizer29_wait = (~main_mon_bussynchronizer29_ping_i);
assign main_mon_bussynchronizer29_ping_i = ((main_mon_bussynchronizer29_starter | main_mon_bussynchronizer29_pong_o) | main_mon_bussynchronizer29_done);
assign main_mon_bussynchronizer29_pong_i = main_mon_bussynchronizer29_ping_o1;
assign main_mon_bussynchronizer29_ping_o0 = (main_mon_bussynchronizer29_ping_toggle_o ^ main_mon_bussynchronizer29_ping_toggle_o_r);
assign main_mon_bussynchronizer29_pong_o = (main_mon_bussynchronizer29_pong_toggle_o ^ main_mon_bussynchronizer29_pong_toggle_o_r);
assign main_mon_bussynchronizer29_done = (main_mon_bussynchronizer29_count == 1'd0);
assign main_mon_bussynchronizer30_wait = (~main_mon_bussynchronizer30_ping_i);
assign main_mon_bussynchronizer30_ping_i = ((main_mon_bussynchronizer30_starter | main_mon_bussynchronizer30_pong_o) | main_mon_bussynchronizer30_done);
assign main_mon_bussynchronizer30_pong_i = main_mon_bussynchronizer30_ping_o1;
assign main_mon_bussynchronizer30_ping_o0 = (main_mon_bussynchronizer30_ping_toggle_o ^ main_mon_bussynchronizer30_ping_toggle_o_r);
assign main_mon_bussynchronizer30_pong_o = (main_mon_bussynchronizer30_pong_toggle_o ^ main_mon_bussynchronizer30_pong_toggle_o_r);
assign main_mon_bussynchronizer30_done = (main_mon_bussynchronizer30_count == 1'd0);
assign main_mon_bussynchronizer31_wait = (~main_mon_bussynchronizer31_ping_i);
assign main_mon_bussynchronizer31_ping_i = ((main_mon_bussynchronizer31_starter | main_mon_bussynchronizer31_pong_o) | main_mon_bussynchronizer31_done);
assign main_mon_bussynchronizer31_pong_i = main_mon_bussynchronizer31_ping_o1;
assign main_mon_bussynchronizer31_ping_o0 = (main_mon_bussynchronizer31_ping_toggle_o ^ main_mon_bussynchronizer31_ping_toggle_o_r);
assign main_mon_bussynchronizer31_pong_o = (main_mon_bussynchronizer31_pong_toggle_o ^ main_mon_bussynchronizer31_pong_toggle_o_r);
assign main_mon_bussynchronizer31_done = (main_mon_bussynchronizer31_count == 1'd0);
assign main_mon_bussynchronizer32_wait = (~main_mon_bussynchronizer32_ping_i);
assign main_mon_bussynchronizer32_ping_i = ((main_mon_bussynchronizer32_starter | main_mon_bussynchronizer32_pong_o) | main_mon_bussynchronizer32_done);
assign main_mon_bussynchronizer32_pong_i = main_mon_bussynchronizer32_ping_o1;
assign main_mon_bussynchronizer32_ping_o0 = (main_mon_bussynchronizer32_ping_toggle_o ^ main_mon_bussynchronizer32_ping_toggle_o_r);
assign main_mon_bussynchronizer32_pong_o = (main_mon_bussynchronizer32_pong_toggle_o ^ main_mon_bussynchronizer32_pong_toggle_o_r);
assign main_mon_bussynchronizer32_done = (main_mon_bussynchronizer32_count == 1'd0);
assign main_mon_bussynchronizer33_wait = (~main_mon_bussynchronizer33_ping_i);
assign main_mon_bussynchronizer33_ping_i = ((main_mon_bussynchronizer33_starter | main_mon_bussynchronizer33_pong_o) | main_mon_bussynchronizer33_done);
assign main_mon_bussynchronizer33_pong_i = main_mon_bussynchronizer33_ping_o1;
assign main_mon_bussynchronizer33_ping_o0 = (main_mon_bussynchronizer33_ping_toggle_o ^ main_mon_bussynchronizer33_ping_toggle_o_r);
assign main_mon_bussynchronizer33_pong_o = (main_mon_bussynchronizer33_pong_toggle_o ^ main_mon_bussynchronizer33_pong_toggle_o_r);
assign main_mon_bussynchronizer33_done = (main_mon_bussynchronizer33_count == 1'd0);
assign main_mon_bussynchronizer34_wait = (~main_mon_bussynchronizer34_ping_i);
assign main_mon_bussynchronizer34_ping_i = ((main_mon_bussynchronizer34_starter | main_mon_bussynchronizer34_pong_o) | main_mon_bussynchronizer34_done);
assign main_mon_bussynchronizer34_pong_i = main_mon_bussynchronizer34_ping_o1;
assign main_mon_bussynchronizer34_ping_o0 = (main_mon_bussynchronizer34_ping_toggle_o ^ main_mon_bussynchronizer34_ping_toggle_o_r);
assign main_mon_bussynchronizer34_pong_o = (main_mon_bussynchronizer34_pong_toggle_o ^ main_mon_bussynchronizer34_pong_toggle_o_r);
assign main_mon_bussynchronizer34_done = (main_mon_bussynchronizer34_count == 1'd0);
assign main_mon_bussynchronizer35_wait = (~main_mon_bussynchronizer35_ping_i);
assign main_mon_bussynchronizer35_ping_i = ((main_mon_bussynchronizer35_starter | main_mon_bussynchronizer35_pong_o) | main_mon_bussynchronizer35_done);
assign main_mon_bussynchronizer35_pong_i = main_mon_bussynchronizer35_ping_o1;
assign main_mon_bussynchronizer35_ping_o0 = (main_mon_bussynchronizer35_ping_toggle_o ^ main_mon_bussynchronizer35_ping_toggle_o_r);
assign main_mon_bussynchronizer35_pong_o = (main_mon_bussynchronizer35_pong_toggle_o ^ main_mon_bussynchronizer35_pong_toggle_o_r);
assign main_mon_bussynchronizer35_done = (main_mon_bussynchronizer35_count == 1'd0);
assign main_mon_bussynchronizer36_wait = (~main_mon_bussynchronizer36_ping_i);
assign main_mon_bussynchronizer36_ping_i = ((main_mon_bussynchronizer36_starter | main_mon_bussynchronizer36_pong_o) | main_mon_bussynchronizer36_done);
assign main_mon_bussynchronizer36_pong_i = main_mon_bussynchronizer36_ping_o1;
assign main_mon_bussynchronizer36_ping_o0 = (main_mon_bussynchronizer36_ping_toggle_o ^ main_mon_bussynchronizer36_ping_toggle_o_r);
assign main_mon_bussynchronizer36_pong_o = (main_mon_bussynchronizer36_pong_toggle_o ^ main_mon_bussynchronizer36_pong_toggle_o_r);
assign main_mon_bussynchronizer36_done = (main_mon_bussynchronizer36_count == 1'd0);
assign main_mon_bussynchronizer37_wait = (~main_mon_bussynchronizer37_ping_i);
assign main_mon_bussynchronizer37_ping_i = ((main_mon_bussynchronizer37_starter | main_mon_bussynchronizer37_pong_o) | main_mon_bussynchronizer37_done);
assign main_mon_bussynchronizer37_pong_i = main_mon_bussynchronizer37_ping_o1;
assign main_mon_bussynchronizer37_ping_o0 = (main_mon_bussynchronizer37_ping_toggle_o ^ main_mon_bussynchronizer37_ping_toggle_o_r);
assign main_mon_bussynchronizer37_pong_o = (main_mon_bussynchronizer37_pong_toggle_o ^ main_mon_bussynchronizer37_pong_toggle_o_r);
assign main_mon_bussynchronizer37_done = (main_mon_bussynchronizer37_count == 1'd0);
assign main_mon_bussynchronizer38_wait = (~main_mon_bussynchronizer38_ping_i);
assign main_mon_bussynchronizer38_ping_i = ((main_mon_bussynchronizer38_starter | main_mon_bussynchronizer38_pong_o) | main_mon_bussynchronizer38_done);
assign main_mon_bussynchronizer38_pong_i = main_mon_bussynchronizer38_ping_o1;
assign main_mon_bussynchronizer38_ping_o0 = (main_mon_bussynchronizer38_ping_toggle_o ^ main_mon_bussynchronizer38_ping_toggle_o_r);
assign main_mon_bussynchronizer38_pong_o = (main_mon_bussynchronizer38_pong_toggle_o ^ main_mon_bussynchronizer38_pong_toggle_o_r);
assign main_mon_bussynchronizer38_done = (main_mon_bussynchronizer38_count == 1'd0);
assign main_inj_value_w = builder_comb_rhs_array_muxed16;
assign main_rtio_analyzer_fifo_sink_stb = main_rtio_analyzer_message_encoder_source_stb;
assign main_rtio_analyzer_message_encoder_source_ack = main_rtio_analyzer_fifo_sink_ack;
assign main_rtio_analyzer_fifo_sink_eop = main_rtio_analyzer_message_encoder_source_eop;
assign main_rtio_analyzer_fifo_sink_payload_data = main_rtio_analyzer_message_encoder_source_payload_data;
assign main_rtio_analyzer_converter_sink_stb = main_rtio_analyzer_fifo_source_stb;
assign main_rtio_analyzer_fifo_source_ack = main_rtio_analyzer_converter_sink_ack;
assign main_rtio_analyzer_converter_sink_eop = main_rtio_analyzer_fifo_source_eop;
assign main_rtio_analyzer_converter_sink_payload_data = main_rtio_analyzer_fifo_source_payload_data;
assign main_rtio_analyzer_dma_sink_stb = main_rtio_analyzer_converter_source_stb;
assign main_rtio_analyzer_converter_source_ack = main_rtio_analyzer_dma_sink_ack;
assign main_rtio_analyzer_dma_sink_eop = main_rtio_analyzer_converter_source_eop;
assign main_rtio_analyzer_dma_sink_payload_data = main_rtio_analyzer_converter_source_payload_data;
assign main_rtio_analyzer_dma_sink_payload_valid_token_count = main_rtio_analyzer_converter_source_payload_valid_token_count;

// synthesis translate_off
reg dummy_d_168;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_read_done <= 1'd0;
	main_rtio_analyzer_message_encoder_read_overflow <= 1'd0;
	if ((main_rtio_analyzer_message_encoder_read_wait_event_r & (~main_rtio_core_cri_i_status[2]))) begin
		if ((~main_rtio_core_cri_i_status[0])) begin
			main_rtio_analyzer_message_encoder_read_done <= 1'd1;
		end
		if (main_rtio_core_cri_i_status[1]) begin
			main_rtio_analyzer_message_encoder_read_overflow <= 1'd1;
		end
	end
// synthesis translate_off
	dummy_d_168 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_input_output_channel = main_rtio_core_cri_chan_sel;
assign main_rtio_analyzer_message_encoder_input_output_address_padding = main_rtio_core_cri_o_address;
assign main_rtio_analyzer_message_encoder_input_output_rtio_counter = main_full_ts_sys;

// synthesis translate_off
reg dummy_d_169;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_input_output_message_type <= 2'd0;
	main_rtio_analyzer_message_encoder_input_output_timestamp <= 64'd0;
	main_rtio_analyzer_message_encoder_input_output_data <= 64'd0;
	if ((main_rtio_core_cri_cmd == 1'd1)) begin
		main_rtio_analyzer_message_encoder_input_output_message_type <= 1'd0;
		main_rtio_analyzer_message_encoder_input_output_timestamp <= main_rtio_core_cri_o_timestamp;
		main_rtio_analyzer_message_encoder_input_output_data <= main_rtio_core_cri_o_data;
	end else begin
		main_rtio_analyzer_message_encoder_input_output_message_type <= 1'd1;
		main_rtio_analyzer_message_encoder_input_output_timestamp <= main_rtio_core_cri_i_timestamp;
		main_rtio_analyzer_message_encoder_input_output_data <= main_rtio_core_cri_i_data;
	end
// synthesis translate_off
	dummy_d_169 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_input_output_stb = ((main_rtio_core_cri_cmd == 1'd1) | main_rtio_analyzer_message_encoder_read_done);
assign main_rtio_analyzer_message_encoder_exception_message_type = 2'd2;
assign main_rtio_analyzer_message_encoder_exception_channel = main_rtio_core_cri_chan_sel;
assign main_rtio_analyzer_message_encoder_exception_rtio_counter = main_full_ts_sys;

// synthesis translate_off
reg dummy_d_170;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_message_encoder_exception_stb <= 1'd0;
	main_rtio_analyzer_message_encoder_exception_exception_type <= 8'd0;
	if ((main_rtio_analyzer_message_encoder_just_written & main_rtio_core_cri_o_status[1])) begin
		main_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_rtio_analyzer_message_encoder_exception_exception_type <= 5'd20;
	end
	if (main_rtio_analyzer_message_encoder_read_overflow) begin
		main_rtio_analyzer_message_encoder_exception_stb <= 1'd1;
		main_rtio_analyzer_message_encoder_exception_exception_type <= 6'd33;
	end
// synthesis translate_off
	dummy_d_170 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_message_encoder_stopped_message_type = 2'd3;
assign main_rtio_analyzer_message_encoder_stopped_rtio_counter = main_full_ts_sys;
assign main_rtio_analyzer_fifo_syncfifo_din = {main_rtio_analyzer_fifo_fifo_in_eop, main_rtio_analyzer_fifo_fifo_in_payload_data};
assign {main_rtio_analyzer_fifo_fifo_out_eop, main_rtio_analyzer_fifo_fifo_out_payload_data} = main_rtio_analyzer_fifo_syncfifo_dout;
assign main_rtio_analyzer_fifo_sink_ack = main_rtio_analyzer_fifo_syncfifo_writable;
assign main_rtio_analyzer_fifo_syncfifo_we = main_rtio_analyzer_fifo_sink_stb;
assign main_rtio_analyzer_fifo_fifo_in_eop = main_rtio_analyzer_fifo_sink_eop;
assign main_rtio_analyzer_fifo_fifo_in_payload_data = main_rtio_analyzer_fifo_sink_payload_data;
assign main_rtio_analyzer_fifo_source_stb = main_rtio_analyzer_fifo_readable;
assign main_rtio_analyzer_fifo_source_eop = main_rtio_analyzer_fifo_fifo_out_eop;
assign main_rtio_analyzer_fifo_source_payload_data = main_rtio_analyzer_fifo_fifo_out_payload_data;
assign main_rtio_analyzer_fifo_re = main_rtio_analyzer_fifo_source_ack;
assign main_rtio_analyzer_fifo_syncfifo_re = (main_rtio_analyzer_fifo_syncfifo_readable & ((~main_rtio_analyzer_fifo_readable) | main_rtio_analyzer_fifo_re));
assign main_rtio_analyzer_fifo_level1 = (main_rtio_analyzer_fifo_level0 + main_rtio_analyzer_fifo_readable);

// synthesis translate_off
reg dummy_d_171;
// synthesis translate_on
always @(*) begin
	main_rtio_analyzer_fifo_wrport_adr <= 7'd0;
	if (main_rtio_analyzer_fifo_replace) begin
		main_rtio_analyzer_fifo_wrport_adr <= (main_rtio_analyzer_fifo_produce - 1'd1);
	end else begin
		main_rtio_analyzer_fifo_wrport_adr <= main_rtio_analyzer_fifo_produce;
	end
// synthesis translate_off
	dummy_d_171 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_fifo_wrport_dat_w = main_rtio_analyzer_fifo_syncfifo_din;
assign main_rtio_analyzer_fifo_wrport_we = (main_rtio_analyzer_fifo_syncfifo_we & (main_rtio_analyzer_fifo_syncfifo_writable | main_rtio_analyzer_fifo_replace));
assign main_rtio_analyzer_fifo_do_read = (main_rtio_analyzer_fifo_syncfifo_readable & main_rtio_analyzer_fifo_syncfifo_re);
assign main_rtio_analyzer_fifo_rdport_adr = main_rtio_analyzer_fifo_consume;
assign main_rtio_analyzer_fifo_syncfifo_dout = main_rtio_analyzer_fifo_rdport_dat_r;
assign main_rtio_analyzer_fifo_rdport_re = main_rtio_analyzer_fifo_do_read;
assign main_rtio_analyzer_fifo_syncfifo_writable = (main_rtio_analyzer_fifo_level0 != 8'd128);
assign main_rtio_analyzer_fifo_syncfifo_readable = (main_rtio_analyzer_fifo_level0 != 1'd0);
assign main_rtio_analyzer_converter_sink_ack = ((~main_rtio_analyzer_converter_strobe_all) | main_rtio_analyzer_converter_source_ack);
assign main_rtio_analyzer_converter_source_stb = main_rtio_analyzer_converter_strobe_all;
assign main_rtio_analyzer_converter_load_part = (main_rtio_analyzer_converter_sink_stb & main_rtio_analyzer_converter_sink_ack);
assign main_interface1_bus_cyc = main_rtio_analyzer_dma_sink_stb;
assign main_interface1_bus_stb = main_rtio_analyzer_dma_sink_stb;
assign main_rtio_analyzer_dma_sink_ack = main_interface1_bus_ack;
assign main_interface1_bus_we = 1'd1;
assign main_interface1_bus_dat_w = main_rtio_analyzer_dma_sink_payload_data;

// synthesis translate_off
reg dummy_d_172;
// synthesis translate_on
always @(*) begin
	main_interface1_bus_sel <= 64'd0;
	main_interface1_bus_sel[0] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[1] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[2] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[3] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[4] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[5] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[6] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[7] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[8] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[9] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[10] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[11] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[12] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[13] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[14] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[15] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[16] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[17] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[18] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[19] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[20] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[21] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[22] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[23] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[24] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[25] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[26] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[27] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[28] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[29] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[30] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[31] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd0);
	main_interface1_bus_sel[32] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[33] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[34] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[35] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[36] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[37] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[38] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[39] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[40] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[41] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[42] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[43] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[44] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[45] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[46] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[47] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[48] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[49] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[50] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[51] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[52] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[53] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[54] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[55] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[56] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[57] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[58] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[59] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[60] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[61] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[62] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
	main_interface1_bus_sel[63] <= (main_rtio_analyzer_dma_sink_payload_valid_token_count >= 1'd1);
// synthesis translate_off
	dummy_d_172 <= dummy_s;
// synthesis translate_on
end
assign main_rtio_analyzer_dma_status = (main_rtio_analyzer_dma_message_count <<< 3'd5);
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr = builder_comb_rhs_array_muxed46;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_w = builder_comb_rhs_array_muxed47;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_sel = builder_comb_rhs_array_muxed48;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cyc = builder_comb_rhs_array_muxed49;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_stb = builder_comb_rhs_array_muxed50;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_we = builder_comb_rhs_array_muxed51;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_cti = builder_comb_rhs_array_muxed52;
assign main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_bte = builder_comb_rhs_array_muxed53;
assign main_nist_clock_nist_clock_wb_sdram_dat_r = main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r;
assign main_kernel_cpu_wb_sdram_dat_r = main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_dat_r;
assign main_nist_clock_nist_clock_wb_sdram_ack = (main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_kernel_cpu_wb_sdram_ack = (main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_ack & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign main_nist_clock_nist_clock_wb_sdram_err = (main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd0));
assign main_kernel_cpu_wb_sdram_err = (main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_err & (builder_sdram_cpulevel_arbiter_grant == 1'd1));
assign builder_sdram_cpulevel_arbiter_request = {(main_kernel_cpu_wb_sdram_cyc & (~main_kernel_cpu_wb_sdram_ack)), (main_nist_clock_nist_clock_wb_sdram_cyc & (~main_nist_clock_nist_clock_wb_sdram_ack))};
assign main_nist_clock_nist_clock_sdram_controller_bus_adr = builder_comb_rhs_array_muxed54;
assign main_nist_clock_nist_clock_sdram_controller_bus_dat_w = builder_comb_rhs_array_muxed55;
assign main_nist_clock_nist_clock_sdram_controller_bus_sel = builder_comb_rhs_array_muxed56;
assign main_nist_clock_nist_clock_sdram_controller_bus_cyc = builder_comb_rhs_array_muxed57;
assign main_nist_clock_nist_clock_sdram_controller_bus_stb = builder_comb_rhs_array_muxed58;
assign main_nist_clock_nist_clock_sdram_controller_bus_we = builder_comb_rhs_array_muxed59;
assign main_nist_clock_nist_clock_sdram_controller_bus_cti = builder_comb_rhs_array_muxed60;
assign main_nist_clock_nist_clock_sdram_controller_bus_bte = builder_comb_rhs_array_muxed61;
assign main_nist_clock_nist_clock_bridge_if_bus_dat_r = main_nist_clock_nist_clock_sdram_controller_bus_dat_r;
assign main_interface0_bus_dat_r = main_nist_clock_nist_clock_sdram_controller_bus_dat_r;
assign main_interface1_bus_dat_r = main_nist_clock_nist_clock_sdram_controller_bus_dat_r;
assign main_nist_clock_nist_clock_bridge_if_bus_ack = (main_nist_clock_nist_clock_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_interface0_bus_ack = (main_nist_clock_nist_clock_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_interface1_bus_ack = (main_nist_clock_nist_clock_sdram_controller_bus_ack & (builder_sdram_native_arbiter_grant == 2'd2));
assign main_nist_clock_nist_clock_bridge_if_bus_err = (main_nist_clock_nist_clock_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd0));
assign main_interface0_bus_err = (main_nist_clock_nist_clock_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 1'd1));
assign main_interface1_bus_err = (main_nist_clock_nist_clock_sdram_controller_bus_err & (builder_sdram_native_arbiter_grant == 2'd2));
assign builder_sdram_native_arbiter_request = {(main_interface1_bus_cyc & (~main_interface1_bus_ack)), (main_interface0_bus_cyc & (~main_interface0_bus_ack)), (main_nist_clock_nist_clock_bridge_if_bus_cyc & (~main_nist_clock_nist_clock_bridge_if_bus_ack))};
assign builder_nist_clock_shared_adr = builder_comb_rhs_array_muxed62;
assign builder_nist_clock_shared_dat_w = builder_comb_rhs_array_muxed63;
assign builder_nist_clock_shared_sel = builder_comb_rhs_array_muxed64;
assign builder_nist_clock_shared_cyc = builder_comb_rhs_array_muxed65;
assign builder_nist_clock_shared_stb = builder_comb_rhs_array_muxed66;
assign builder_nist_clock_shared_we = builder_comb_rhs_array_muxed67;
assign builder_nist_clock_shared_cti = builder_comb_rhs_array_muxed68;
assign builder_nist_clock_shared_bte = builder_comb_rhs_array_muxed69;
assign main_nist_clock_nist_clock_ibus_dat_r = builder_nist_clock_shared_dat_r;
assign main_nist_clock_nist_clock_tmpu_dat_r = builder_nist_clock_shared_dat_r;
assign main_nist_clock_nist_clock_ibus_ack = (builder_nist_clock_shared_ack & (builder_nist_clock_grant == 1'd0));
assign main_nist_clock_nist_clock_tmpu_ack = (builder_nist_clock_shared_ack & (builder_nist_clock_grant == 1'd1));
assign main_nist_clock_nist_clock_ibus_err = (builder_nist_clock_shared_err & (builder_nist_clock_grant == 1'd0));
assign main_nist_clock_nist_clock_tmpu_err = (builder_nist_clock_shared_err & (builder_nist_clock_grant == 1'd1));
assign builder_nist_clock_request = {(main_nist_clock_nist_clock_tmpu_cyc & (~main_nist_clock_nist_clock_tmpu_ack)), (main_nist_clock_nist_clock_ibus_cyc & (~main_nist_clock_nist_clock_ibus_ack))};

// synthesis translate_off
reg dummy_d_173;
// synthesis translate_on
always @(*) begin
	builder_nist_clock_slave_sel <= 6'd0;
	builder_nist_clock_slave_sel[0] <= (((1'd1 & (~builder_nist_clock_shared_adr[27])) & (~builder_nist_clock_shared_adr[28])) & builder_nist_clock_shared_adr[26]);
	builder_nist_clock_slave_sel[1] <= (((1'd1 & (~builder_nist_clock_shared_adr[26])) & builder_nist_clock_shared_adr[27]) & builder_nist_clock_shared_adr[28]);
	builder_nist_clock_slave_sel[2] <= ((1'd1 & (~builder_nist_clock_shared_adr[27])) & builder_nist_clock_shared_adr[28]);
	builder_nist_clock_slave_sel[3] <= (((1'd1 & (~builder_nist_clock_shared_adr[26])) & (~builder_nist_clock_shared_adr[27])) & (~builder_nist_clock_shared_adr[28]));
	builder_nist_clock_slave_sel[4] <= ((1'd1 & (~builder_nist_clock_shared_adr[28])) & builder_nist_clock_shared_adr[27]);
	builder_nist_clock_slave_sel[5] <= (((1'd1 & builder_nist_clock_shared_adr[26]) & builder_nist_clock_shared_adr[27]) & builder_nist_clock_shared_adr[28]);
// synthesis translate_off
	dummy_d_173 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_sram_bus_adr = builder_nist_clock_shared_adr;
assign main_nist_clock_nist_clock_sram_bus_dat_w = builder_nist_clock_shared_dat_w;
assign main_nist_clock_nist_clock_sram_bus_sel = builder_nist_clock_shared_sel;
assign main_nist_clock_nist_clock_sram_bus_stb = builder_nist_clock_shared_stb;
assign main_nist_clock_nist_clock_sram_bus_we = builder_nist_clock_shared_we;
assign main_nist_clock_nist_clock_sram_bus_cti = builder_nist_clock_shared_cti;
assign main_nist_clock_nist_clock_sram_bus_bte = builder_nist_clock_shared_bte;
assign main_nist_clock_nist_clock_bus_wishbone_adr = builder_nist_clock_shared_adr;
assign main_nist_clock_nist_clock_bus_wishbone_dat_w = builder_nist_clock_shared_dat_w;
assign main_nist_clock_nist_clock_bus_wishbone_sel = builder_nist_clock_shared_sel;
assign main_nist_clock_nist_clock_bus_wishbone_stb = builder_nist_clock_shared_stb;
assign main_nist_clock_nist_clock_bus_wishbone_we = builder_nist_clock_shared_we;
assign main_nist_clock_nist_clock_bus_wishbone_cti = builder_nist_clock_shared_cti;
assign main_nist_clock_nist_clock_bus_wishbone_bte = builder_nist_clock_shared_bte;
assign main_nist_clock_nist_clock_wb_sdram_adr = builder_nist_clock_shared_adr;
assign main_nist_clock_nist_clock_wb_sdram_dat_w = builder_nist_clock_shared_dat_w;
assign main_nist_clock_nist_clock_wb_sdram_sel = builder_nist_clock_shared_sel;
assign main_nist_clock_nist_clock_wb_sdram_stb = builder_nist_clock_shared_stb;
assign main_nist_clock_nist_clock_wb_sdram_we = builder_nist_clock_shared_we;
assign main_nist_clock_nist_clock_wb_sdram_cti = builder_nist_clock_shared_cti;
assign main_nist_clock_nist_clock_wb_sdram_bte = builder_nist_clock_shared_bte;
assign main_nist_clock_spiflash_bus_adr = builder_nist_clock_shared_adr;
assign main_nist_clock_spiflash_bus_dat_w = builder_nist_clock_shared_dat_w;
assign main_nist_clock_spiflash_bus_sel = builder_nist_clock_shared_sel;
assign main_nist_clock_spiflash_bus_stb = builder_nist_clock_shared_stb;
assign main_nist_clock_spiflash_bus_we = builder_nist_clock_shared_we;
assign main_nist_clock_spiflash_bus_cti = builder_nist_clock_shared_cti;
assign main_nist_clock_spiflash_bus_bte = builder_nist_clock_shared_bte;
assign main_bus_adr = builder_nist_clock_shared_adr;
assign main_bus_dat_w = builder_nist_clock_shared_dat_w;
assign main_bus_sel = builder_nist_clock_shared_sel;
assign main_bus_stb = builder_nist_clock_shared_stb;
assign main_bus_we = builder_nist_clock_shared_we;
assign main_bus_cti = builder_nist_clock_shared_cti;
assign main_bus_bte = builder_nist_clock_shared_bte;
assign main_mailbox_i1_adr = builder_nist_clock_shared_adr;
assign main_mailbox_i1_dat_w = builder_nist_clock_shared_dat_w;
assign main_mailbox_i1_sel = builder_nist_clock_shared_sel;
assign main_mailbox_i1_stb = builder_nist_clock_shared_stb;
assign main_mailbox_i1_we = builder_nist_clock_shared_we;
assign main_mailbox_i1_cti = builder_nist_clock_shared_cti;
assign main_mailbox_i1_bte = builder_nist_clock_shared_bte;
assign main_nist_clock_nist_clock_sram_bus_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[0]);
assign main_nist_clock_nist_clock_bus_wishbone_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[1]);
assign main_nist_clock_nist_clock_wb_sdram_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[2]);
assign main_nist_clock_spiflash_bus_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[3]);
assign main_bus_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[4]);
assign main_mailbox_i1_cyc = (builder_nist_clock_shared_cyc & builder_nist_clock_slave_sel[5]);
assign builder_nist_clock_shared_ack = (((((main_nist_clock_nist_clock_sram_bus_ack | main_nist_clock_nist_clock_bus_wishbone_ack) | main_nist_clock_nist_clock_wb_sdram_ack) | main_nist_clock_spiflash_bus_ack) | main_bus_ack) | main_mailbox_i1_ack);
assign builder_nist_clock_shared_err = (((((main_nist_clock_nist_clock_sram_bus_err | main_nist_clock_nist_clock_bus_wishbone_err) | main_nist_clock_nist_clock_wb_sdram_err) | main_nist_clock_spiflash_bus_err) | main_bus_err) | main_mailbox_i1_err);
assign builder_nist_clock_shared_dat_r = (((((({32{builder_nist_clock_slave_sel_r[0]}} & main_nist_clock_nist_clock_sram_bus_dat_r) | ({32{builder_nist_clock_slave_sel_r[1]}} & main_nist_clock_nist_clock_bus_wishbone_dat_r)) | ({32{builder_nist_clock_slave_sel_r[2]}} & main_nist_clock_nist_clock_wb_sdram_dat_r)) | ({32{builder_nist_clock_slave_sel_r[3]}} & main_nist_clock_spiflash_bus_dat_r)) | ({32{builder_nist_clock_slave_sel_r[4]}} & main_bus_dat_r)) | ({32{builder_nist_clock_slave_sel_r[5]}} & main_mailbox_i1_dat_r));
assign builder_nist_clock_csrbank0_sel = (builder_nist_clock_interface0_bank_bus_adr[13:9] == 3'd7);
assign builder_nist_clock_csrbank0_wlevel_en0_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank0_wlevel_en0_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 1'd0));
assign main_nist_clock_ddrphy_wlevel_strobe_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_wlevel_strobe_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 1'd1));
assign builder_nist_clock_csrbank0_dly_sel0_r = builder_nist_clock_interface0_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank0_dly_sel0_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 2'd2));
assign main_nist_clock_ddrphy_rdly_dq_rst_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_rdly_dq_rst_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 2'd3));
assign main_nist_clock_ddrphy_rdly_dq_inc_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_rdly_dq_inc_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 3'd4));
assign main_nist_clock_ddrphy_rdly_dq_bitslip_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_rdly_dq_bitslip_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 3'd5));
assign main_nist_clock_ddrphy_wdly_dq_rst_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_wdly_dq_rst_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 3'd6));
assign main_nist_clock_ddrphy_wdly_dq_inc_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_wdly_dq_inc_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 3'd7));
assign main_nist_clock_ddrphy_wdly_dqs_rst_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_wdly_dqs_rst_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 4'd8));
assign main_nist_clock_ddrphy_wdly_dqs_inc_r = builder_nist_clock_interface0_bank_bus_dat_w[0];
assign main_nist_clock_ddrphy_wdly_dqs_inc_re = ((builder_nist_clock_csrbank0_sel & builder_nist_clock_interface0_bank_bus_we) & (builder_nist_clock_interface0_bank_bus_adr[3:0] == 4'd9));
assign main_nist_clock_ddrphy_wlevel_en_storage = main_nist_clock_ddrphy_wlevel_en_storage_full;
assign builder_nist_clock_csrbank0_wlevel_en0_w = main_nist_clock_ddrphy_wlevel_en_storage_full;
assign main_nist_clock_ddrphy_dly_sel_storage = main_nist_clock_ddrphy_dly_sel_storage_full[7:0];
assign builder_nist_clock_csrbank0_dly_sel0_w = main_nist_clock_ddrphy_dly_sel_storage_full[7:0];
assign builder_nist_clock_csrbank1_sel = (builder_nist_clock_interface1_bank_bus_adr[13:9] == 3'd5);
assign builder_nist_clock_csrbank1_control0_r = builder_nist_clock_interface1_bank_bus_dat_w[3:0];
assign builder_nist_clock_csrbank1_control0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 1'd0));
assign builder_nist_clock_csrbank1_pi0_command0_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi0_command0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 1'd1));
assign main_nist_clock_nist_clock_phaseinjector0_command_issue_r = builder_nist_clock_interface1_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_phaseinjector0_command_issue_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 2'd2));
assign builder_nist_clock_csrbank1_pi0_address1_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi0_address1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 2'd3));
assign builder_nist_clock_csrbank1_pi0_address0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_address0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 3'd4));
assign builder_nist_clock_csrbank1_pi0_baddress0_r = builder_nist_clock_interface1_bank_bus_dat_w[2:0];
assign builder_nist_clock_csrbank1_pi0_baddress0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 3'd5));
assign builder_nist_clock_csrbank1_pi0_wrdata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 3'd6));
assign builder_nist_clock_csrbank1_pi0_wrdata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 3'd7));
assign builder_nist_clock_csrbank1_pi0_wrdata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd8));
assign builder_nist_clock_csrbank1_pi0_wrdata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd9));
assign builder_nist_clock_csrbank1_pi0_wrdata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd10));
assign builder_nist_clock_csrbank1_pi0_wrdata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd11));
assign builder_nist_clock_csrbank1_pi0_wrdata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd12));
assign builder_nist_clock_csrbank1_pi0_wrdata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd13));
assign builder_nist_clock_csrbank1_pi0_wrdata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd14));
assign builder_nist_clock_csrbank1_pi0_wrdata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 4'd15));
assign builder_nist_clock_csrbank1_pi0_wrdata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd16));
assign builder_nist_clock_csrbank1_pi0_wrdata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd17));
assign builder_nist_clock_csrbank1_pi0_wrdata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd18));
assign builder_nist_clock_csrbank1_pi0_wrdata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd19));
assign builder_nist_clock_csrbank1_pi0_wrdata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd20));
assign builder_nist_clock_csrbank1_pi0_wrdata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_wrdata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd21));
assign builder_nist_clock_csrbank1_pi0_rddata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd22));
assign builder_nist_clock_csrbank1_pi0_rddata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd23));
assign builder_nist_clock_csrbank1_pi0_rddata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd24));
assign builder_nist_clock_csrbank1_pi0_rddata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd25));
assign builder_nist_clock_csrbank1_pi0_rddata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd26));
assign builder_nist_clock_csrbank1_pi0_rddata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd27));
assign builder_nist_clock_csrbank1_pi0_rddata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd28));
assign builder_nist_clock_csrbank1_pi0_rddata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd29));
assign builder_nist_clock_csrbank1_pi0_rddata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd30));
assign builder_nist_clock_csrbank1_pi0_rddata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 5'd31));
assign builder_nist_clock_csrbank1_pi0_rddata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd32));
assign builder_nist_clock_csrbank1_pi0_rddata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd33));
assign builder_nist_clock_csrbank1_pi0_rddata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd34));
assign builder_nist_clock_csrbank1_pi0_rddata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd35));
assign builder_nist_clock_csrbank1_pi0_rddata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd36));
assign builder_nist_clock_csrbank1_pi0_rddata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd37));
assign builder_nist_clock_csrbank1_pi1_command0_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi1_command0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd38));
assign main_nist_clock_nist_clock_phaseinjector1_command_issue_r = builder_nist_clock_interface1_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_phaseinjector1_command_issue_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd39));
assign builder_nist_clock_csrbank1_pi1_address1_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi1_address1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd40));
assign builder_nist_clock_csrbank1_pi1_address0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_address0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd41));
assign builder_nist_clock_csrbank1_pi1_baddress0_r = builder_nist_clock_interface1_bank_bus_dat_w[2:0];
assign builder_nist_clock_csrbank1_pi1_baddress0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd42));
assign builder_nist_clock_csrbank1_pi1_wrdata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd43));
assign builder_nist_clock_csrbank1_pi1_wrdata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd44));
assign builder_nist_clock_csrbank1_pi1_wrdata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd45));
assign builder_nist_clock_csrbank1_pi1_wrdata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd46));
assign builder_nist_clock_csrbank1_pi1_wrdata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd47));
assign builder_nist_clock_csrbank1_pi1_wrdata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd48));
assign builder_nist_clock_csrbank1_pi1_wrdata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd49));
assign builder_nist_clock_csrbank1_pi1_wrdata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd50));
assign builder_nist_clock_csrbank1_pi1_wrdata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd51));
assign builder_nist_clock_csrbank1_pi1_wrdata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd52));
assign builder_nist_clock_csrbank1_pi1_wrdata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd53));
assign builder_nist_clock_csrbank1_pi1_wrdata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd54));
assign builder_nist_clock_csrbank1_pi1_wrdata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd55));
assign builder_nist_clock_csrbank1_pi1_wrdata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd56));
assign builder_nist_clock_csrbank1_pi1_wrdata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd57));
assign builder_nist_clock_csrbank1_pi1_wrdata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_wrdata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd58));
assign builder_nist_clock_csrbank1_pi1_rddata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd59));
assign builder_nist_clock_csrbank1_pi1_rddata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd60));
assign builder_nist_clock_csrbank1_pi1_rddata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd61));
assign builder_nist_clock_csrbank1_pi1_rddata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd62));
assign builder_nist_clock_csrbank1_pi1_rddata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 6'd63));
assign builder_nist_clock_csrbank1_pi1_rddata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd64));
assign builder_nist_clock_csrbank1_pi1_rddata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd65));
assign builder_nist_clock_csrbank1_pi1_rddata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd66));
assign builder_nist_clock_csrbank1_pi1_rddata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd67));
assign builder_nist_clock_csrbank1_pi1_rddata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd68));
assign builder_nist_clock_csrbank1_pi1_rddata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd69));
assign builder_nist_clock_csrbank1_pi1_rddata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd70));
assign builder_nist_clock_csrbank1_pi1_rddata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd71));
assign builder_nist_clock_csrbank1_pi1_rddata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd72));
assign builder_nist_clock_csrbank1_pi1_rddata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd73));
assign builder_nist_clock_csrbank1_pi1_rddata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd74));
assign builder_nist_clock_csrbank1_pi2_command0_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi2_command0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd75));
assign main_nist_clock_nist_clock_phaseinjector2_command_issue_r = builder_nist_clock_interface1_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_phaseinjector2_command_issue_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd76));
assign builder_nist_clock_csrbank1_pi2_address1_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi2_address1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd77));
assign builder_nist_clock_csrbank1_pi2_address0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_address0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd78));
assign builder_nist_clock_csrbank1_pi2_baddress0_r = builder_nist_clock_interface1_bank_bus_dat_w[2:0];
assign builder_nist_clock_csrbank1_pi2_baddress0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd79));
assign builder_nist_clock_csrbank1_pi2_wrdata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd80));
assign builder_nist_clock_csrbank1_pi2_wrdata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd81));
assign builder_nist_clock_csrbank1_pi2_wrdata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd82));
assign builder_nist_clock_csrbank1_pi2_wrdata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd83));
assign builder_nist_clock_csrbank1_pi2_wrdata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd84));
assign builder_nist_clock_csrbank1_pi2_wrdata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd85));
assign builder_nist_clock_csrbank1_pi2_wrdata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd86));
assign builder_nist_clock_csrbank1_pi2_wrdata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd87));
assign builder_nist_clock_csrbank1_pi2_wrdata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd88));
assign builder_nist_clock_csrbank1_pi2_wrdata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd89));
assign builder_nist_clock_csrbank1_pi2_wrdata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd90));
assign builder_nist_clock_csrbank1_pi2_wrdata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd91));
assign builder_nist_clock_csrbank1_pi2_wrdata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd92));
assign builder_nist_clock_csrbank1_pi2_wrdata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd93));
assign builder_nist_clock_csrbank1_pi2_wrdata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd94));
assign builder_nist_clock_csrbank1_pi2_wrdata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_wrdata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd95));
assign builder_nist_clock_csrbank1_pi2_rddata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd96));
assign builder_nist_clock_csrbank1_pi2_rddata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd97));
assign builder_nist_clock_csrbank1_pi2_rddata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd98));
assign builder_nist_clock_csrbank1_pi2_rddata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd99));
assign builder_nist_clock_csrbank1_pi2_rddata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd100));
assign builder_nist_clock_csrbank1_pi2_rddata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd101));
assign builder_nist_clock_csrbank1_pi2_rddata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd102));
assign builder_nist_clock_csrbank1_pi2_rddata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd103));
assign builder_nist_clock_csrbank1_pi2_rddata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd104));
assign builder_nist_clock_csrbank1_pi2_rddata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd105));
assign builder_nist_clock_csrbank1_pi2_rddata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd106));
assign builder_nist_clock_csrbank1_pi2_rddata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd107));
assign builder_nist_clock_csrbank1_pi2_rddata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd108));
assign builder_nist_clock_csrbank1_pi2_rddata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd109));
assign builder_nist_clock_csrbank1_pi2_rddata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd110));
assign builder_nist_clock_csrbank1_pi2_rddata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd111));
assign builder_nist_clock_csrbank1_pi3_command0_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi3_command0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd112));
assign main_nist_clock_nist_clock_phaseinjector3_command_issue_r = builder_nist_clock_interface1_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_phaseinjector3_command_issue_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd113));
assign builder_nist_clock_csrbank1_pi3_address1_r = builder_nist_clock_interface1_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank1_pi3_address1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd114));
assign builder_nist_clock_csrbank1_pi3_address0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_address0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd115));
assign builder_nist_clock_csrbank1_pi3_baddress0_r = builder_nist_clock_interface1_bank_bus_dat_w[2:0];
assign builder_nist_clock_csrbank1_pi3_baddress0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd116));
assign builder_nist_clock_csrbank1_pi3_wrdata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd117));
assign builder_nist_clock_csrbank1_pi3_wrdata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd118));
assign builder_nist_clock_csrbank1_pi3_wrdata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd119));
assign builder_nist_clock_csrbank1_pi3_wrdata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd120));
assign builder_nist_clock_csrbank1_pi3_wrdata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd121));
assign builder_nist_clock_csrbank1_pi3_wrdata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd122));
assign builder_nist_clock_csrbank1_pi3_wrdata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd123));
assign builder_nist_clock_csrbank1_pi3_wrdata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd124));
assign builder_nist_clock_csrbank1_pi3_wrdata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd125));
assign builder_nist_clock_csrbank1_pi3_wrdata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd126));
assign builder_nist_clock_csrbank1_pi3_wrdata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 7'd127));
assign builder_nist_clock_csrbank1_pi3_wrdata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd128));
assign builder_nist_clock_csrbank1_pi3_wrdata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd129));
assign builder_nist_clock_csrbank1_pi3_wrdata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd130));
assign builder_nist_clock_csrbank1_pi3_wrdata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd131));
assign builder_nist_clock_csrbank1_pi3_wrdata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_wrdata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd132));
assign builder_nist_clock_csrbank1_pi3_rddata15_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata15_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd133));
assign builder_nist_clock_csrbank1_pi3_rddata14_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata14_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd134));
assign builder_nist_clock_csrbank1_pi3_rddata13_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata13_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd135));
assign builder_nist_clock_csrbank1_pi3_rddata12_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata12_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd136));
assign builder_nist_clock_csrbank1_pi3_rddata11_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata11_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd137));
assign builder_nist_clock_csrbank1_pi3_rddata10_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata10_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd138));
assign builder_nist_clock_csrbank1_pi3_rddata9_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata9_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd139));
assign builder_nist_clock_csrbank1_pi3_rddata8_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata8_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd140));
assign builder_nist_clock_csrbank1_pi3_rddata7_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata7_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd141));
assign builder_nist_clock_csrbank1_pi3_rddata6_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata6_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd142));
assign builder_nist_clock_csrbank1_pi3_rddata5_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata5_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd143));
assign builder_nist_clock_csrbank1_pi3_rddata4_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata4_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd144));
assign builder_nist_clock_csrbank1_pi3_rddata3_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata3_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd145));
assign builder_nist_clock_csrbank1_pi3_rddata2_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata2_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd146));
assign builder_nist_clock_csrbank1_pi3_rddata1_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata1_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd147));
assign builder_nist_clock_csrbank1_pi3_rddata0_r = builder_nist_clock_interface1_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata0_re = ((builder_nist_clock_csrbank1_sel & builder_nist_clock_interface1_bank_bus_we) & (builder_nist_clock_interface1_bank_bus_adr[7:0] == 8'd148));
assign main_nist_clock_nist_clock_storage = main_nist_clock_nist_clock_storage_full[3:0];
assign builder_nist_clock_csrbank1_control0_w = main_nist_clock_nist_clock_storage_full[3:0];
assign main_nist_clock_nist_clock_phaseinjector0_command_storage = main_nist_clock_nist_clock_phaseinjector0_command_storage_full[5:0];
assign builder_nist_clock_csrbank1_pi0_command0_w = main_nist_clock_nist_clock_phaseinjector0_command_storage_full[5:0];
assign main_nist_clock_nist_clock_phaseinjector0_address_storage = main_nist_clock_nist_clock_phaseinjector0_address_storage_full[13:0];
assign builder_nist_clock_csrbank1_pi0_address1_w = main_nist_clock_nist_clock_phaseinjector0_address_storage_full[13:8];
assign builder_nist_clock_csrbank1_pi0_address0_w = main_nist_clock_nist_clock_phaseinjector0_address_storage_full[7:0];
assign main_nist_clock_nist_clock_phaseinjector0_baddress_storage = main_nist_clock_nist_clock_phaseinjector0_baddress_storage_full[2:0];
assign builder_nist_clock_csrbank1_pi0_baddress0_w = main_nist_clock_nist_clock_phaseinjector0_baddress_storage_full[2:0];
assign main_nist_clock_nist_clock_phaseinjector0_wrdata_storage = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[127:0];
assign builder_nist_clock_csrbank1_pi0_wrdata15_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[127:120];
assign builder_nist_clock_csrbank1_pi0_wrdata14_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[119:112];
assign builder_nist_clock_csrbank1_pi0_wrdata13_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[111:104];
assign builder_nist_clock_csrbank1_pi0_wrdata12_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[103:96];
assign builder_nist_clock_csrbank1_pi0_wrdata11_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[95:88];
assign builder_nist_clock_csrbank1_pi0_wrdata10_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[87:80];
assign builder_nist_clock_csrbank1_pi0_wrdata9_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[79:72];
assign builder_nist_clock_csrbank1_pi0_wrdata8_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[71:64];
assign builder_nist_clock_csrbank1_pi0_wrdata7_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[63:56];
assign builder_nist_clock_csrbank1_pi0_wrdata6_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[55:48];
assign builder_nist_clock_csrbank1_pi0_wrdata5_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[47:40];
assign builder_nist_clock_csrbank1_pi0_wrdata4_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[39:32];
assign builder_nist_clock_csrbank1_pi0_wrdata3_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[31:24];
assign builder_nist_clock_csrbank1_pi0_wrdata2_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[23:16];
assign builder_nist_clock_csrbank1_pi0_wrdata1_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[15:8];
assign builder_nist_clock_csrbank1_pi0_wrdata0_w = main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[7:0];
assign builder_nist_clock_csrbank1_pi0_rddata15_w = main_nist_clock_nist_clock_phaseinjector0_status[127:120];
assign builder_nist_clock_csrbank1_pi0_rddata14_w = main_nist_clock_nist_clock_phaseinjector0_status[119:112];
assign builder_nist_clock_csrbank1_pi0_rddata13_w = main_nist_clock_nist_clock_phaseinjector0_status[111:104];
assign builder_nist_clock_csrbank1_pi0_rddata12_w = main_nist_clock_nist_clock_phaseinjector0_status[103:96];
assign builder_nist_clock_csrbank1_pi0_rddata11_w = main_nist_clock_nist_clock_phaseinjector0_status[95:88];
assign builder_nist_clock_csrbank1_pi0_rddata10_w = main_nist_clock_nist_clock_phaseinjector0_status[87:80];
assign builder_nist_clock_csrbank1_pi0_rddata9_w = main_nist_clock_nist_clock_phaseinjector0_status[79:72];
assign builder_nist_clock_csrbank1_pi0_rddata8_w = main_nist_clock_nist_clock_phaseinjector0_status[71:64];
assign builder_nist_clock_csrbank1_pi0_rddata7_w = main_nist_clock_nist_clock_phaseinjector0_status[63:56];
assign builder_nist_clock_csrbank1_pi0_rddata6_w = main_nist_clock_nist_clock_phaseinjector0_status[55:48];
assign builder_nist_clock_csrbank1_pi0_rddata5_w = main_nist_clock_nist_clock_phaseinjector0_status[47:40];
assign builder_nist_clock_csrbank1_pi0_rddata4_w = main_nist_clock_nist_clock_phaseinjector0_status[39:32];
assign builder_nist_clock_csrbank1_pi0_rddata3_w = main_nist_clock_nist_clock_phaseinjector0_status[31:24];
assign builder_nist_clock_csrbank1_pi0_rddata2_w = main_nist_clock_nist_clock_phaseinjector0_status[23:16];
assign builder_nist_clock_csrbank1_pi0_rddata1_w = main_nist_clock_nist_clock_phaseinjector0_status[15:8];
assign builder_nist_clock_csrbank1_pi0_rddata0_w = main_nist_clock_nist_clock_phaseinjector0_status[7:0];
assign main_nist_clock_nist_clock_phaseinjector1_command_storage = main_nist_clock_nist_clock_phaseinjector1_command_storage_full[5:0];
assign builder_nist_clock_csrbank1_pi1_command0_w = main_nist_clock_nist_clock_phaseinjector1_command_storage_full[5:0];
assign main_nist_clock_nist_clock_phaseinjector1_address_storage = main_nist_clock_nist_clock_phaseinjector1_address_storage_full[13:0];
assign builder_nist_clock_csrbank1_pi1_address1_w = main_nist_clock_nist_clock_phaseinjector1_address_storage_full[13:8];
assign builder_nist_clock_csrbank1_pi1_address0_w = main_nist_clock_nist_clock_phaseinjector1_address_storage_full[7:0];
assign main_nist_clock_nist_clock_phaseinjector1_baddress_storage = main_nist_clock_nist_clock_phaseinjector1_baddress_storage_full[2:0];
assign builder_nist_clock_csrbank1_pi1_baddress0_w = main_nist_clock_nist_clock_phaseinjector1_baddress_storage_full[2:0];
assign main_nist_clock_nist_clock_phaseinjector1_wrdata_storage = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[127:0];
assign builder_nist_clock_csrbank1_pi1_wrdata15_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[127:120];
assign builder_nist_clock_csrbank1_pi1_wrdata14_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[119:112];
assign builder_nist_clock_csrbank1_pi1_wrdata13_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[111:104];
assign builder_nist_clock_csrbank1_pi1_wrdata12_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[103:96];
assign builder_nist_clock_csrbank1_pi1_wrdata11_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[95:88];
assign builder_nist_clock_csrbank1_pi1_wrdata10_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[87:80];
assign builder_nist_clock_csrbank1_pi1_wrdata9_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[79:72];
assign builder_nist_clock_csrbank1_pi1_wrdata8_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[71:64];
assign builder_nist_clock_csrbank1_pi1_wrdata7_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[63:56];
assign builder_nist_clock_csrbank1_pi1_wrdata6_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[55:48];
assign builder_nist_clock_csrbank1_pi1_wrdata5_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[47:40];
assign builder_nist_clock_csrbank1_pi1_wrdata4_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[39:32];
assign builder_nist_clock_csrbank1_pi1_wrdata3_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[31:24];
assign builder_nist_clock_csrbank1_pi1_wrdata2_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[23:16];
assign builder_nist_clock_csrbank1_pi1_wrdata1_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[15:8];
assign builder_nist_clock_csrbank1_pi1_wrdata0_w = main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[7:0];
assign builder_nist_clock_csrbank1_pi1_rddata15_w = main_nist_clock_nist_clock_phaseinjector1_status[127:120];
assign builder_nist_clock_csrbank1_pi1_rddata14_w = main_nist_clock_nist_clock_phaseinjector1_status[119:112];
assign builder_nist_clock_csrbank1_pi1_rddata13_w = main_nist_clock_nist_clock_phaseinjector1_status[111:104];
assign builder_nist_clock_csrbank1_pi1_rddata12_w = main_nist_clock_nist_clock_phaseinjector1_status[103:96];
assign builder_nist_clock_csrbank1_pi1_rddata11_w = main_nist_clock_nist_clock_phaseinjector1_status[95:88];
assign builder_nist_clock_csrbank1_pi1_rddata10_w = main_nist_clock_nist_clock_phaseinjector1_status[87:80];
assign builder_nist_clock_csrbank1_pi1_rddata9_w = main_nist_clock_nist_clock_phaseinjector1_status[79:72];
assign builder_nist_clock_csrbank1_pi1_rddata8_w = main_nist_clock_nist_clock_phaseinjector1_status[71:64];
assign builder_nist_clock_csrbank1_pi1_rddata7_w = main_nist_clock_nist_clock_phaseinjector1_status[63:56];
assign builder_nist_clock_csrbank1_pi1_rddata6_w = main_nist_clock_nist_clock_phaseinjector1_status[55:48];
assign builder_nist_clock_csrbank1_pi1_rddata5_w = main_nist_clock_nist_clock_phaseinjector1_status[47:40];
assign builder_nist_clock_csrbank1_pi1_rddata4_w = main_nist_clock_nist_clock_phaseinjector1_status[39:32];
assign builder_nist_clock_csrbank1_pi1_rddata3_w = main_nist_clock_nist_clock_phaseinjector1_status[31:24];
assign builder_nist_clock_csrbank1_pi1_rddata2_w = main_nist_clock_nist_clock_phaseinjector1_status[23:16];
assign builder_nist_clock_csrbank1_pi1_rddata1_w = main_nist_clock_nist_clock_phaseinjector1_status[15:8];
assign builder_nist_clock_csrbank1_pi1_rddata0_w = main_nist_clock_nist_clock_phaseinjector1_status[7:0];
assign main_nist_clock_nist_clock_phaseinjector2_command_storage = main_nist_clock_nist_clock_phaseinjector2_command_storage_full[5:0];
assign builder_nist_clock_csrbank1_pi2_command0_w = main_nist_clock_nist_clock_phaseinjector2_command_storage_full[5:0];
assign main_nist_clock_nist_clock_phaseinjector2_address_storage = main_nist_clock_nist_clock_phaseinjector2_address_storage_full[13:0];
assign builder_nist_clock_csrbank1_pi2_address1_w = main_nist_clock_nist_clock_phaseinjector2_address_storage_full[13:8];
assign builder_nist_clock_csrbank1_pi2_address0_w = main_nist_clock_nist_clock_phaseinjector2_address_storage_full[7:0];
assign main_nist_clock_nist_clock_phaseinjector2_baddress_storage = main_nist_clock_nist_clock_phaseinjector2_baddress_storage_full[2:0];
assign builder_nist_clock_csrbank1_pi2_baddress0_w = main_nist_clock_nist_clock_phaseinjector2_baddress_storage_full[2:0];
assign main_nist_clock_nist_clock_phaseinjector2_wrdata_storage = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[127:0];
assign builder_nist_clock_csrbank1_pi2_wrdata15_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[127:120];
assign builder_nist_clock_csrbank1_pi2_wrdata14_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[119:112];
assign builder_nist_clock_csrbank1_pi2_wrdata13_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[111:104];
assign builder_nist_clock_csrbank1_pi2_wrdata12_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[103:96];
assign builder_nist_clock_csrbank1_pi2_wrdata11_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[95:88];
assign builder_nist_clock_csrbank1_pi2_wrdata10_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[87:80];
assign builder_nist_clock_csrbank1_pi2_wrdata9_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[79:72];
assign builder_nist_clock_csrbank1_pi2_wrdata8_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[71:64];
assign builder_nist_clock_csrbank1_pi2_wrdata7_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[63:56];
assign builder_nist_clock_csrbank1_pi2_wrdata6_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[55:48];
assign builder_nist_clock_csrbank1_pi2_wrdata5_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[47:40];
assign builder_nist_clock_csrbank1_pi2_wrdata4_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[39:32];
assign builder_nist_clock_csrbank1_pi2_wrdata3_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[31:24];
assign builder_nist_clock_csrbank1_pi2_wrdata2_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[23:16];
assign builder_nist_clock_csrbank1_pi2_wrdata1_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[15:8];
assign builder_nist_clock_csrbank1_pi2_wrdata0_w = main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[7:0];
assign builder_nist_clock_csrbank1_pi2_rddata15_w = main_nist_clock_nist_clock_phaseinjector2_status[127:120];
assign builder_nist_clock_csrbank1_pi2_rddata14_w = main_nist_clock_nist_clock_phaseinjector2_status[119:112];
assign builder_nist_clock_csrbank1_pi2_rddata13_w = main_nist_clock_nist_clock_phaseinjector2_status[111:104];
assign builder_nist_clock_csrbank1_pi2_rddata12_w = main_nist_clock_nist_clock_phaseinjector2_status[103:96];
assign builder_nist_clock_csrbank1_pi2_rddata11_w = main_nist_clock_nist_clock_phaseinjector2_status[95:88];
assign builder_nist_clock_csrbank1_pi2_rddata10_w = main_nist_clock_nist_clock_phaseinjector2_status[87:80];
assign builder_nist_clock_csrbank1_pi2_rddata9_w = main_nist_clock_nist_clock_phaseinjector2_status[79:72];
assign builder_nist_clock_csrbank1_pi2_rddata8_w = main_nist_clock_nist_clock_phaseinjector2_status[71:64];
assign builder_nist_clock_csrbank1_pi2_rddata7_w = main_nist_clock_nist_clock_phaseinjector2_status[63:56];
assign builder_nist_clock_csrbank1_pi2_rddata6_w = main_nist_clock_nist_clock_phaseinjector2_status[55:48];
assign builder_nist_clock_csrbank1_pi2_rddata5_w = main_nist_clock_nist_clock_phaseinjector2_status[47:40];
assign builder_nist_clock_csrbank1_pi2_rddata4_w = main_nist_clock_nist_clock_phaseinjector2_status[39:32];
assign builder_nist_clock_csrbank1_pi2_rddata3_w = main_nist_clock_nist_clock_phaseinjector2_status[31:24];
assign builder_nist_clock_csrbank1_pi2_rddata2_w = main_nist_clock_nist_clock_phaseinjector2_status[23:16];
assign builder_nist_clock_csrbank1_pi2_rddata1_w = main_nist_clock_nist_clock_phaseinjector2_status[15:8];
assign builder_nist_clock_csrbank1_pi2_rddata0_w = main_nist_clock_nist_clock_phaseinjector2_status[7:0];
assign main_nist_clock_nist_clock_phaseinjector3_command_storage = main_nist_clock_nist_clock_phaseinjector3_command_storage_full[5:0];
assign builder_nist_clock_csrbank1_pi3_command0_w = main_nist_clock_nist_clock_phaseinjector3_command_storage_full[5:0];
assign main_nist_clock_nist_clock_phaseinjector3_address_storage = main_nist_clock_nist_clock_phaseinjector3_address_storage_full[13:0];
assign builder_nist_clock_csrbank1_pi3_address1_w = main_nist_clock_nist_clock_phaseinjector3_address_storage_full[13:8];
assign builder_nist_clock_csrbank1_pi3_address0_w = main_nist_clock_nist_clock_phaseinjector3_address_storage_full[7:0];
assign main_nist_clock_nist_clock_phaseinjector3_baddress_storage = main_nist_clock_nist_clock_phaseinjector3_baddress_storage_full[2:0];
assign builder_nist_clock_csrbank1_pi3_baddress0_w = main_nist_clock_nist_clock_phaseinjector3_baddress_storage_full[2:0];
assign main_nist_clock_nist_clock_phaseinjector3_wrdata_storage = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[127:0];
assign builder_nist_clock_csrbank1_pi3_wrdata15_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[127:120];
assign builder_nist_clock_csrbank1_pi3_wrdata14_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[119:112];
assign builder_nist_clock_csrbank1_pi3_wrdata13_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[111:104];
assign builder_nist_clock_csrbank1_pi3_wrdata12_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[103:96];
assign builder_nist_clock_csrbank1_pi3_wrdata11_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[95:88];
assign builder_nist_clock_csrbank1_pi3_wrdata10_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[87:80];
assign builder_nist_clock_csrbank1_pi3_wrdata9_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[79:72];
assign builder_nist_clock_csrbank1_pi3_wrdata8_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[71:64];
assign builder_nist_clock_csrbank1_pi3_wrdata7_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[63:56];
assign builder_nist_clock_csrbank1_pi3_wrdata6_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[55:48];
assign builder_nist_clock_csrbank1_pi3_wrdata5_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[47:40];
assign builder_nist_clock_csrbank1_pi3_wrdata4_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[39:32];
assign builder_nist_clock_csrbank1_pi3_wrdata3_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[31:24];
assign builder_nist_clock_csrbank1_pi3_wrdata2_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[23:16];
assign builder_nist_clock_csrbank1_pi3_wrdata1_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[15:8];
assign builder_nist_clock_csrbank1_pi3_wrdata0_w = main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[7:0];
assign builder_nist_clock_csrbank1_pi3_rddata15_w = main_nist_clock_nist_clock_phaseinjector3_status[127:120];
assign builder_nist_clock_csrbank1_pi3_rddata14_w = main_nist_clock_nist_clock_phaseinjector3_status[119:112];
assign builder_nist_clock_csrbank1_pi3_rddata13_w = main_nist_clock_nist_clock_phaseinjector3_status[111:104];
assign builder_nist_clock_csrbank1_pi3_rddata12_w = main_nist_clock_nist_clock_phaseinjector3_status[103:96];
assign builder_nist_clock_csrbank1_pi3_rddata11_w = main_nist_clock_nist_clock_phaseinjector3_status[95:88];
assign builder_nist_clock_csrbank1_pi3_rddata10_w = main_nist_clock_nist_clock_phaseinjector3_status[87:80];
assign builder_nist_clock_csrbank1_pi3_rddata9_w = main_nist_clock_nist_clock_phaseinjector3_status[79:72];
assign builder_nist_clock_csrbank1_pi3_rddata8_w = main_nist_clock_nist_clock_phaseinjector3_status[71:64];
assign builder_nist_clock_csrbank1_pi3_rddata7_w = main_nist_clock_nist_clock_phaseinjector3_status[63:56];
assign builder_nist_clock_csrbank1_pi3_rddata6_w = main_nist_clock_nist_clock_phaseinjector3_status[55:48];
assign builder_nist_clock_csrbank1_pi3_rddata5_w = main_nist_clock_nist_clock_phaseinjector3_status[47:40];
assign builder_nist_clock_csrbank1_pi3_rddata4_w = main_nist_clock_nist_clock_phaseinjector3_status[39:32];
assign builder_nist_clock_csrbank1_pi3_rddata3_w = main_nist_clock_nist_clock_phaseinjector3_status[31:24];
assign builder_nist_clock_csrbank1_pi3_rddata2_w = main_nist_clock_nist_clock_phaseinjector3_status[23:16];
assign builder_nist_clock_csrbank1_pi3_rddata1_w = main_nist_clock_nist_clock_phaseinjector3_status[15:8];
assign builder_nist_clock_csrbank1_pi3_rddata0_w = main_nist_clock_nist_clock_phaseinjector3_status[7:0];
assign builder_nist_clock_csrbank2_sel = (builder_nist_clock_interface2_bank_bus_adr[13:9] == 4'd10);
assign builder_nist_clock_csrbank2_sram_writer_slot_r = builder_nist_clock_interface2_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank2_sram_writer_slot_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 1'd0));
assign builder_nist_clock_csrbank2_sram_writer_length3_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_length3_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 1'd1));
assign builder_nist_clock_csrbank2_sram_writer_length2_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_length2_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 2'd2));
assign builder_nist_clock_csrbank2_sram_writer_length1_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_length1_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 2'd3));
assign builder_nist_clock_csrbank2_sram_writer_length0_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_length0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 3'd4));
assign builder_nist_clock_csrbank2_sram_writer_errors3_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_errors3_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 3'd5));
assign builder_nist_clock_csrbank2_sram_writer_errors2_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_errors2_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 3'd6));
assign builder_nist_clock_csrbank2_sram_writer_errors1_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_errors1_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 3'd7));
assign builder_nist_clock_csrbank2_sram_writer_errors0_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_writer_errors0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd8));
assign main_writer_status_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign main_writer_status_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd9));
assign main_writer_pending_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign main_writer_pending_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd10));
assign builder_nist_clock_csrbank2_sram_writer_ev_enable0_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank2_sram_writer_ev_enable0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd11));
assign main_reader_start_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign main_reader_start_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd12));
assign builder_nist_clock_csrbank2_sram_reader_ready_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank2_sram_reader_ready_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd13));
assign builder_nist_clock_csrbank2_sram_reader_slot0_r = builder_nist_clock_interface2_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank2_sram_reader_slot0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd14));
assign builder_nist_clock_csrbank2_sram_reader_length1_r = builder_nist_clock_interface2_bank_bus_dat_w[2:0];
assign builder_nist_clock_csrbank2_sram_reader_length1_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 4'd15));
assign builder_nist_clock_csrbank2_sram_reader_length0_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_sram_reader_length0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd16));
assign main_reader_eventmanager_status_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign main_reader_eventmanager_status_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd17));
assign main_reader_eventmanager_pending_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign main_reader_eventmanager_pending_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd18));
assign builder_nist_clock_csrbank2_sram_reader_ev_enable0_r = builder_nist_clock_interface2_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank2_sram_reader_ev_enable0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd19));
assign builder_nist_clock_csrbank2_preamble_errors3_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_preamble_errors3_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd20));
assign builder_nist_clock_csrbank2_preamble_errors2_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_preamble_errors2_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd21));
assign builder_nist_clock_csrbank2_preamble_errors1_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_preamble_errors1_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd22));
assign builder_nist_clock_csrbank2_preamble_errors0_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_preamble_errors0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd23));
assign builder_nist_clock_csrbank2_crc_errors3_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_crc_errors3_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd24));
assign builder_nist_clock_csrbank2_crc_errors2_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_crc_errors2_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd25));
assign builder_nist_clock_csrbank2_crc_errors1_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_crc_errors1_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd26));
assign builder_nist_clock_csrbank2_crc_errors0_r = builder_nist_clock_interface2_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank2_crc_errors0_re = ((builder_nist_clock_csrbank2_sel & builder_nist_clock_interface2_bank_bus_we) & (builder_nist_clock_interface2_bank_bus_adr[4:0] == 5'd27));
assign builder_nist_clock_csrbank2_sram_writer_slot_w = main_writer_slot_status[1:0];
assign builder_nist_clock_csrbank2_sram_writer_length3_w = main_writer_length_status[31:24];
assign builder_nist_clock_csrbank2_sram_writer_length2_w = main_writer_length_status[23:16];
assign builder_nist_clock_csrbank2_sram_writer_length1_w = main_writer_length_status[15:8];
assign builder_nist_clock_csrbank2_sram_writer_length0_w = main_writer_length_status[7:0];
assign builder_nist_clock_csrbank2_sram_writer_errors3_w = main_writer_errors_status[31:24];
assign builder_nist_clock_csrbank2_sram_writer_errors2_w = main_writer_errors_status[23:16];
assign builder_nist_clock_csrbank2_sram_writer_errors1_w = main_writer_errors_status[15:8];
assign builder_nist_clock_csrbank2_sram_writer_errors0_w = main_writer_errors_status[7:0];
assign main_writer_storage = main_writer_storage_full;
assign builder_nist_clock_csrbank2_sram_writer_ev_enable0_w = main_writer_storage_full;
assign builder_nist_clock_csrbank2_sram_reader_ready_w = main_reader_ready_status;
assign main_reader_slot_storage = main_reader_slot_storage_full[1:0];
assign builder_nist_clock_csrbank2_sram_reader_slot0_w = main_reader_slot_storage_full[1:0];
assign main_reader_length_storage = main_reader_length_storage_full[10:0];
assign builder_nist_clock_csrbank2_sram_reader_length1_w = main_reader_length_storage_full[10:8];
assign builder_nist_clock_csrbank2_sram_reader_length0_w = main_reader_length_storage_full[7:0];
assign main_reader_eventmanager_storage = main_reader_eventmanager_storage_full;
assign builder_nist_clock_csrbank2_sram_reader_ev_enable0_w = main_reader_eventmanager_storage_full;
assign builder_nist_clock_csrbank2_preamble_errors3_w = main_preamble_errors_status[31:24];
assign builder_nist_clock_csrbank2_preamble_errors2_w = main_preamble_errors_status[23:16];
assign builder_nist_clock_csrbank2_preamble_errors1_w = main_preamble_errors_status[15:8];
assign builder_nist_clock_csrbank2_preamble_errors0_w = main_preamble_errors_status[7:0];
assign builder_nist_clock_csrbank2_crc_errors3_w = main_crc_errors_status[31:24];
assign builder_nist_clock_csrbank2_crc_errors2_w = main_crc_errors_status[23:16];
assign builder_nist_clock_csrbank2_crc_errors1_w = main_crc_errors_status[15:8];
assign builder_nist_clock_csrbank2_crc_errors0_w = main_crc_errors_status[7:0];
assign builder_nist_clock_csrbank3_sel = (builder_nist_clock_interface3_bank_bus_adr[13:9] == 4'd9);
assign builder_nist_clock_csrbank3_mode_detection_mode_r = builder_nist_clock_interface3_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank3_mode_detection_mode_re = ((builder_nist_clock_csrbank3_sel & builder_nist_clock_interface3_bank_bus_we) & (builder_nist_clock_interface3_bank_bus_adr[0] == 1'd0));
assign builder_nist_clock_csrbank3_crg_reset0_r = builder_nist_clock_interface3_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank3_crg_reset0_re = ((builder_nist_clock_csrbank3_sel & builder_nist_clock_interface3_bank_bus_we) & (builder_nist_clock_interface3_bank_bus_adr[0] == 1'd1));
assign builder_nist_clock_csrbank3_mode_detection_mode_w = main_ethphy_mode_status;
assign main_ethphy_storage = main_ethphy_storage_full;
assign builder_nist_clock_csrbank3_crg_reset0_w = main_ethphy_storage_full;
assign builder_nist_clock_csrbank4_sel = (builder_nist_clock_interface4_bank_bus_adr[13:9] == 4'd14);
assign builder_nist_clock_csrbank4_in_r = builder_nist_clock_interface4_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank4_in_re = ((builder_nist_clock_csrbank4_sel & builder_nist_clock_interface4_bank_bus_we) & (builder_nist_clock_interface4_bank_bus_adr[1:0] == 1'd0));
assign builder_nist_clock_csrbank4_out0_r = builder_nist_clock_interface4_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank4_out0_re = ((builder_nist_clock_csrbank4_sel & builder_nist_clock_interface4_bank_bus_we) & (builder_nist_clock_interface4_bank_bus_adr[1:0] == 1'd1));
assign builder_nist_clock_csrbank4_oe0_r = builder_nist_clock_interface4_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank4_oe0_re = ((builder_nist_clock_csrbank4_sel & builder_nist_clock_interface4_bank_bus_we) & (builder_nist_clock_interface4_bank_bus_adr[1:0] == 2'd2));
assign builder_nist_clock_csrbank4_in_w = main_i2c_status0[1:0];
assign main_i2c_out_storage = main_i2c_out_storage_full[1:0];
assign builder_nist_clock_csrbank4_out0_w = main_i2c_out_storage_full[1:0];
assign main_i2c_oe_storage = main_i2c_oe_storage_full[1:0];
assign builder_nist_clock_csrbank4_oe0_w = main_i2c_oe_storage_full[1:0];
assign builder_nist_clock_csrbank5_sel = (builder_nist_clock_interface5_bank_bus_adr[13:9] == 2'd2);
assign builder_nist_clock_csrbank5_address0_r = builder_nist_clock_interface5_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank5_address0_re = ((builder_nist_clock_csrbank5_sel & builder_nist_clock_interface5_bank_bus_we) & (builder_nist_clock_interface5_bank_bus_adr[0] == 1'd0));
assign builder_nist_clock_csrbank5_data_r = builder_nist_clock_interface5_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank5_data_re = ((builder_nist_clock_csrbank5_sel & builder_nist_clock_interface5_bank_bus_we) & (builder_nist_clock_interface5_bank_bus_adr[0] == 1'd1));
assign main_add_identifier_storage = main_add_identifier_storage_full[7:0];
assign builder_nist_clock_csrbank5_address0_w = main_add_identifier_storage_full[7:0];
assign builder_nist_clock_csrbank5_data_w = main_add_identifier_status[7:0];
assign builder_nist_clock_csrbank6_sel = (builder_nist_clock_interface6_bank_bus_adr[13:9] == 4'd11);
assign builder_nist_clock_csrbank6_reset0_r = builder_nist_clock_interface6_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank6_reset0_re = ((builder_nist_clock_csrbank6_sel & builder_nist_clock_interface6_bank_bus_we) & (builder_nist_clock_interface6_bank_bus_adr[0] == 1'd0));
assign main_kernel_cpu_storage = main_kernel_cpu_storage_full;
assign builder_nist_clock_csrbank6_reset0_w = main_kernel_cpu_storage_full;
assign builder_nist_clock_csrbank7_sel = (builder_nist_clock_interface7_bank_bus_adr[13:9] == 4'd13);
assign builder_nist_clock_csrbank7_out0_r = builder_nist_clock_interface7_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank7_out0_re = ((builder_nist_clock_csrbank7_sel & builder_nist_clock_interface7_bank_bus_we) & (builder_nist_clock_interface7_bank_bus_adr[0] == 1'd0));
assign main_leds_storage = main_leds_storage_full[1:0];
assign builder_nist_clock_csrbank7_out0_w = main_leds_storage_full[1:0];
assign builder_nist_clock_csrbank8_sel = (builder_nist_clock_interface8_bank_bus_adr[13:9] == 5'd18);
assign builder_nist_clock_csrbank8_enable0_r = builder_nist_clock_interface8_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank8_enable0_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 1'd0));
assign builder_nist_clock_csrbank8_busy_r = builder_nist_clock_interface8_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank8_busy_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 1'd1));
assign builder_nist_clock_csrbank8_message_encoder_overflow_r = builder_nist_clock_interface8_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank8_message_encoder_overflow_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 2'd2));
assign main_rtio_analyzer_message_encoder_overflow_reset_r = builder_nist_clock_interface8_bank_bus_dat_w[0];
assign main_rtio_analyzer_message_encoder_overflow_reset_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 2'd3));
assign main_rtio_analyzer_dma_reset_r = builder_nist_clock_interface8_bank_bus_dat_w[0];
assign main_rtio_analyzer_dma_reset_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 3'd4));
assign builder_nist_clock_csrbank8_dma_base_address4_r = builder_nist_clock_interface8_bank_bus_dat_w[3:0];
assign builder_nist_clock_csrbank8_dma_base_address4_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 3'd5));
assign builder_nist_clock_csrbank8_dma_base_address3_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_base_address3_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 3'd6));
assign builder_nist_clock_csrbank8_dma_base_address2_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_base_address2_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 3'd7));
assign builder_nist_clock_csrbank8_dma_base_address1_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_base_address1_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd8));
assign builder_nist_clock_csrbank8_dma_base_address0_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_base_address0_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd9));
assign builder_nist_clock_csrbank8_dma_last_address4_r = builder_nist_clock_interface8_bank_bus_dat_w[3:0];
assign builder_nist_clock_csrbank8_dma_last_address4_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd10));
assign builder_nist_clock_csrbank8_dma_last_address3_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_last_address3_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd11));
assign builder_nist_clock_csrbank8_dma_last_address2_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_last_address2_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd12));
assign builder_nist_clock_csrbank8_dma_last_address1_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_last_address1_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd13));
assign builder_nist_clock_csrbank8_dma_last_address0_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_last_address0_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd14));
assign builder_nist_clock_csrbank8_dma_byte_count7_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count7_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 4'd15));
assign builder_nist_clock_csrbank8_dma_byte_count6_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count6_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd16));
assign builder_nist_clock_csrbank8_dma_byte_count5_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count5_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd17));
assign builder_nist_clock_csrbank8_dma_byte_count4_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count4_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd18));
assign builder_nist_clock_csrbank8_dma_byte_count3_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count3_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd19));
assign builder_nist_clock_csrbank8_dma_byte_count2_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count2_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd20));
assign builder_nist_clock_csrbank8_dma_byte_count1_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count1_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd21));
assign builder_nist_clock_csrbank8_dma_byte_count0_r = builder_nist_clock_interface8_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank8_dma_byte_count0_re = ((builder_nist_clock_csrbank8_sel & builder_nist_clock_interface8_bank_bus_we) & (builder_nist_clock_interface8_bank_bus_adr[4:0] == 5'd22));
assign main_rtio_analyzer_enable_storage = main_rtio_analyzer_enable_storage_full;
assign builder_nist_clock_csrbank8_enable0_w = main_rtio_analyzer_enable_storage_full;
assign builder_nist_clock_csrbank8_busy_w = main_rtio_analyzer_busy_status;
assign builder_nist_clock_csrbank8_message_encoder_overflow_w = main_rtio_analyzer_message_encoder_status;
assign main_rtio_analyzer_dma_base_address_storage = main_rtio_analyzer_dma_base_address_storage_full[35:6];
assign builder_nist_clock_csrbank8_dma_base_address4_w = main_rtio_analyzer_dma_base_address_storage_full[35:32];
assign builder_nist_clock_csrbank8_dma_base_address3_w = main_rtio_analyzer_dma_base_address_storage_full[31:24];
assign builder_nist_clock_csrbank8_dma_base_address2_w = main_rtio_analyzer_dma_base_address_storage_full[23:16];
assign builder_nist_clock_csrbank8_dma_base_address1_w = main_rtio_analyzer_dma_base_address_storage_full[15:8];
assign builder_nist_clock_csrbank8_dma_base_address0_w = {main_rtio_analyzer_dma_base_address_storage_full[7:6], {2{1'd0}}};
assign main_rtio_analyzer_dma_last_address_storage = main_rtio_analyzer_dma_last_address_storage_full[35:6];
assign builder_nist_clock_csrbank8_dma_last_address4_w = main_rtio_analyzer_dma_last_address_storage_full[35:32];
assign builder_nist_clock_csrbank8_dma_last_address3_w = main_rtio_analyzer_dma_last_address_storage_full[31:24];
assign builder_nist_clock_csrbank8_dma_last_address2_w = main_rtio_analyzer_dma_last_address_storage_full[23:16];
assign builder_nist_clock_csrbank8_dma_last_address1_w = main_rtio_analyzer_dma_last_address_storage_full[15:8];
assign builder_nist_clock_csrbank8_dma_last_address0_w = {main_rtio_analyzer_dma_last_address_storage_full[7:6], {2{1'd0}}};
assign builder_nist_clock_csrbank8_dma_byte_count7_w = main_rtio_analyzer_dma_status[63:56];
assign builder_nist_clock_csrbank8_dma_byte_count6_w = main_rtio_analyzer_dma_status[55:48];
assign builder_nist_clock_csrbank8_dma_byte_count5_w = main_rtio_analyzer_dma_status[47:40];
assign builder_nist_clock_csrbank8_dma_byte_count4_w = main_rtio_analyzer_dma_status[39:32];
assign builder_nist_clock_csrbank8_dma_byte_count3_w = main_rtio_analyzer_dma_status[31:24];
assign builder_nist_clock_csrbank8_dma_byte_count2_w = main_rtio_analyzer_dma_status[23:16];
assign builder_nist_clock_csrbank8_dma_byte_count1_w = main_rtio_analyzer_dma_status[15:8];
assign builder_nist_clock_csrbank8_dma_byte_count0_w = main_rtio_analyzer_dma_status[7:0];
assign builder_nist_clock_csrbank9_sel = (builder_nist_clock_interface9_bank_bus_adr[13:9] == 5'd16);
assign main_rtio_core_reset_r = builder_nist_clock_interface9_bank_bus_dat_w[0];
assign main_rtio_core_reset_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 1'd0));
assign main_rtio_core_reset_phy_r = builder_nist_clock_interface9_bank_bus_dat_w[0];
assign main_rtio_core_reset_phy_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 1'd1));
assign main_rtio_core_async_error_r = builder_nist_clock_interface9_bank_bus_dat_w[2:0];
assign main_rtio_core_async_error_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 2'd2));
assign builder_nist_clock_csrbank9_collision_channel1_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_collision_channel1_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 2'd3));
assign builder_nist_clock_csrbank9_collision_channel0_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_collision_channel0_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 3'd4));
assign builder_nist_clock_csrbank9_busy_channel1_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_busy_channel1_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 3'd5));
assign builder_nist_clock_csrbank9_busy_channel0_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_busy_channel0_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 3'd6));
assign builder_nist_clock_csrbank9_sequence_error_channel1_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_sequence_error_channel1_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 3'd7));
assign builder_nist_clock_csrbank9_sequence_error_channel0_r = builder_nist_clock_interface9_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank9_sequence_error_channel0_re = ((builder_nist_clock_csrbank9_sel & builder_nist_clock_interface9_bank_bus_we) & (builder_nist_clock_interface9_bank_bus_adr[3:0] == 4'd8));
assign builder_nist_clock_csrbank9_collision_channel1_w = main_rtio_core_collision_channel_status[15:8];
assign builder_nist_clock_csrbank9_collision_channel0_w = main_rtio_core_collision_channel_status[7:0];
assign builder_nist_clock_csrbank9_busy_channel1_w = main_rtio_core_busy_channel_status[15:8];
assign builder_nist_clock_csrbank9_busy_channel0_w = main_rtio_core_busy_channel_status[7:0];
assign builder_nist_clock_csrbank9_sequence_error_channel1_w = main_rtio_core_sequence_error_channel_status[15:8];
assign builder_nist_clock_csrbank9_sequence_error_channel0_w = main_rtio_core_sequence_error_channel_status[7:0];
assign builder_nist_clock_csrbank10_sel = (builder_nist_clock_interface10_bank_bus_adr[13:9] == 4'd15);
assign builder_nist_clock_csrbank10_clock_sel0_r = builder_nist_clock_interface10_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank10_clock_sel0_re = ((builder_nist_clock_csrbank10_sel & builder_nist_clock_interface10_bank_bus_we) & (builder_nist_clock_interface10_bank_bus_adr[1:0] == 1'd0));
assign builder_nist_clock_csrbank10_pll_reset0_r = builder_nist_clock_interface10_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank10_pll_reset0_re = ((builder_nist_clock_csrbank10_sel & builder_nist_clock_interface10_bank_bus_we) & (builder_nist_clock_interface10_bank_bus_adr[1:0] == 1'd1));
assign builder_nist_clock_csrbank10_pll_locked_r = builder_nist_clock_interface10_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank10_pll_locked_re = ((builder_nist_clock_csrbank10_sel & builder_nist_clock_interface10_bank_bus_we) & (builder_nist_clock_interface10_bank_bus_adr[1:0] == 2'd2));
assign main_rtio_crg_clock_sel_storage = main_rtio_crg_clock_sel_storage_full;
assign builder_nist_clock_csrbank10_clock_sel0_w = main_rtio_crg_clock_sel_storage_full;
assign main_rtio_crg_pll_reset_storage = main_rtio_crg_pll_reset_storage_full;
assign builder_nist_clock_csrbank10_pll_reset0_w = main_rtio_crg_pll_reset_storage_full;
assign builder_nist_clock_csrbank10_pll_locked_w = main_rtio_crg_pll_locked_status;
assign builder_nist_clock_csrbank11_sel = (builder_nist_clock_interface11_bank_bus_adr[13:9] == 5'd17);
assign builder_nist_clock_csrbank11_mon_chan_sel0_r = builder_nist_clock_interface11_bank_bus_dat_w[4:0];
assign builder_nist_clock_csrbank11_mon_chan_sel0_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 1'd0));
assign builder_nist_clock_csrbank11_mon_probe_sel0_r = builder_nist_clock_interface11_bank_bus_dat_w[3:0];
assign builder_nist_clock_csrbank11_mon_probe_sel0_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 1'd1));
assign main_mon_value_update_r = builder_nist_clock_interface11_bank_bus_dat_w[0];
assign main_mon_value_update_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 2'd2));
assign builder_nist_clock_csrbank11_mon_value3_r = builder_nist_clock_interface11_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank11_mon_value3_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 2'd3));
assign builder_nist_clock_csrbank11_mon_value2_r = builder_nist_clock_interface11_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank11_mon_value2_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 3'd4));
assign builder_nist_clock_csrbank11_mon_value1_r = builder_nist_clock_interface11_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank11_mon_value1_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 3'd5));
assign builder_nist_clock_csrbank11_mon_value0_r = builder_nist_clock_interface11_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank11_mon_value0_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 3'd6));
assign builder_nist_clock_csrbank11_inj_chan_sel0_r = builder_nist_clock_interface11_bank_bus_dat_w[4:0];
assign builder_nist_clock_csrbank11_inj_chan_sel0_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 3'd7));
assign builder_nist_clock_csrbank11_inj_override_sel0_r = builder_nist_clock_interface11_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank11_inj_override_sel0_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 4'd8));
assign main_inj_value_r = builder_nist_clock_interface11_bank_bus_dat_w[0];
assign main_inj_value_re = ((builder_nist_clock_csrbank11_sel & builder_nist_clock_interface11_bank_bus_we) & (builder_nist_clock_interface11_bank_bus_adr[3:0] == 4'd9));
assign main_mon_chan_sel_storage = main_mon_chan_sel_storage_full[4:0];
assign builder_nist_clock_csrbank11_mon_chan_sel0_w = main_mon_chan_sel_storage_full[4:0];
assign main_mon_probe_sel_storage = main_mon_probe_sel_storage_full[3:0];
assign builder_nist_clock_csrbank11_mon_probe_sel0_w = main_mon_probe_sel_storage_full[3:0];
assign builder_nist_clock_csrbank11_mon_value3_w = main_mon_status[31:24];
assign builder_nist_clock_csrbank11_mon_value2_w = main_mon_status[23:16];
assign builder_nist_clock_csrbank11_mon_value1_w = main_mon_status[15:8];
assign builder_nist_clock_csrbank11_mon_value0_w = main_mon_status[7:0];
assign main_inj_chan_sel_storage = main_inj_chan_sel_storage_full[4:0];
assign builder_nist_clock_csrbank11_inj_chan_sel0_w = main_inj_chan_sel_storage_full[4:0];
assign main_inj_override_sel_storage = main_inj_override_sel_storage_full[1:0];
assign builder_nist_clock_csrbank11_inj_override_sel0_w = main_inj_override_sel_storage_full[1:0];
assign builder_nist_clock_csrbank12_sel = (builder_nist_clock_interface12_bank_bus_adr[13:9] == 4'd8);
assign builder_nist_clock_csrbank12_bitbang0_r = builder_nist_clock_interface12_bank_bus_dat_w[3:0];
assign builder_nist_clock_csrbank12_bitbang0_re = ((builder_nist_clock_csrbank12_sel & builder_nist_clock_interface12_bank_bus_we) & (builder_nist_clock_interface12_bank_bus_adr[1:0] == 1'd0));
assign builder_nist_clock_csrbank12_miso_r = builder_nist_clock_interface12_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank12_miso_re = ((builder_nist_clock_csrbank12_sel & builder_nist_clock_interface12_bank_bus_we) & (builder_nist_clock_interface12_bank_bus_adr[1:0] == 1'd1));
assign builder_nist_clock_csrbank12_bitbang_en0_r = builder_nist_clock_interface12_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank12_bitbang_en0_re = ((builder_nist_clock_csrbank12_sel & builder_nist_clock_interface12_bank_bus_we) & (builder_nist_clock_interface12_bank_bus_adr[1:0] == 2'd2));
assign main_nist_clock_spiflash_bitbang_storage = main_nist_clock_spiflash_bitbang_storage_full[3:0];
assign builder_nist_clock_csrbank12_bitbang0_w = main_nist_clock_spiflash_bitbang_storage_full[3:0];
assign builder_nist_clock_csrbank12_miso_w = main_nist_clock_spiflash_status;
assign main_nist_clock_spiflash_bitbang_en_storage = main_nist_clock_spiflash_bitbang_en_storage_full;
assign builder_nist_clock_csrbank12_bitbang_en0_w = main_nist_clock_spiflash_bitbang_en_storage_full;
assign builder_nist_clock_csrbank13_sel = (builder_nist_clock_interface13_bank_bus_adr[13:9] == 2'd3);
assign builder_nist_clock_csrbank13_load7_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load7_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 1'd0));
assign builder_nist_clock_csrbank13_load6_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load6_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 1'd1));
assign builder_nist_clock_csrbank13_load5_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load5_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 2'd2));
assign builder_nist_clock_csrbank13_load4_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load4_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 2'd3));
assign builder_nist_clock_csrbank13_load3_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load3_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 3'd4));
assign builder_nist_clock_csrbank13_load2_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load2_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 3'd5));
assign builder_nist_clock_csrbank13_load1_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load1_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 3'd6));
assign builder_nist_clock_csrbank13_load0_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_load0_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 3'd7));
assign builder_nist_clock_csrbank13_reload7_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload7_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd8));
assign builder_nist_clock_csrbank13_reload6_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload6_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd9));
assign builder_nist_clock_csrbank13_reload5_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload5_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd10));
assign builder_nist_clock_csrbank13_reload4_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload4_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd11));
assign builder_nist_clock_csrbank13_reload3_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload3_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd12));
assign builder_nist_clock_csrbank13_reload2_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload2_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd13));
assign builder_nist_clock_csrbank13_reload1_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload1_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd14));
assign builder_nist_clock_csrbank13_reload0_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_reload0_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 4'd15));
assign builder_nist_clock_csrbank13_en0_r = builder_nist_clock_interface13_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank13_en0_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd16));
assign main_nist_clock_nist_clock_timer0_update_value_r = builder_nist_clock_interface13_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_timer0_update_value_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd17));
assign builder_nist_clock_csrbank13_value7_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value7_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd18));
assign builder_nist_clock_csrbank13_value6_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value6_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd19));
assign builder_nist_clock_csrbank13_value5_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value5_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd20));
assign builder_nist_clock_csrbank13_value4_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value4_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd21));
assign builder_nist_clock_csrbank13_value3_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value3_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd22));
assign builder_nist_clock_csrbank13_value2_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value2_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd23));
assign builder_nist_clock_csrbank13_value1_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value1_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd24));
assign builder_nist_clock_csrbank13_value0_r = builder_nist_clock_interface13_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank13_value0_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd25));
assign main_nist_clock_nist_clock_timer0_eventmanager_status_r = builder_nist_clock_interface13_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_timer0_eventmanager_status_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd26));
assign main_nist_clock_nist_clock_timer0_eventmanager_pending_r = builder_nist_clock_interface13_bank_bus_dat_w[0];
assign main_nist_clock_nist_clock_timer0_eventmanager_pending_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd27));
assign builder_nist_clock_csrbank13_ev_enable0_r = builder_nist_clock_interface13_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank13_ev_enable0_re = ((builder_nist_clock_csrbank13_sel & builder_nist_clock_interface13_bank_bus_we) & (builder_nist_clock_interface13_bank_bus_adr[4:0] == 5'd28));
assign main_nist_clock_nist_clock_timer0_load_storage = main_nist_clock_nist_clock_timer0_load_storage_full[63:0];
assign builder_nist_clock_csrbank13_load7_w = main_nist_clock_nist_clock_timer0_load_storage_full[63:56];
assign builder_nist_clock_csrbank13_load6_w = main_nist_clock_nist_clock_timer0_load_storage_full[55:48];
assign builder_nist_clock_csrbank13_load5_w = main_nist_clock_nist_clock_timer0_load_storage_full[47:40];
assign builder_nist_clock_csrbank13_load4_w = main_nist_clock_nist_clock_timer0_load_storage_full[39:32];
assign builder_nist_clock_csrbank13_load3_w = main_nist_clock_nist_clock_timer0_load_storage_full[31:24];
assign builder_nist_clock_csrbank13_load2_w = main_nist_clock_nist_clock_timer0_load_storage_full[23:16];
assign builder_nist_clock_csrbank13_load1_w = main_nist_clock_nist_clock_timer0_load_storage_full[15:8];
assign builder_nist_clock_csrbank13_load0_w = main_nist_clock_nist_clock_timer0_load_storage_full[7:0];
assign main_nist_clock_nist_clock_timer0_reload_storage = main_nist_clock_nist_clock_timer0_reload_storage_full[63:0];
assign builder_nist_clock_csrbank13_reload7_w = main_nist_clock_nist_clock_timer0_reload_storage_full[63:56];
assign builder_nist_clock_csrbank13_reload6_w = main_nist_clock_nist_clock_timer0_reload_storage_full[55:48];
assign builder_nist_clock_csrbank13_reload5_w = main_nist_clock_nist_clock_timer0_reload_storage_full[47:40];
assign builder_nist_clock_csrbank13_reload4_w = main_nist_clock_nist_clock_timer0_reload_storage_full[39:32];
assign builder_nist_clock_csrbank13_reload3_w = main_nist_clock_nist_clock_timer0_reload_storage_full[31:24];
assign builder_nist_clock_csrbank13_reload2_w = main_nist_clock_nist_clock_timer0_reload_storage_full[23:16];
assign builder_nist_clock_csrbank13_reload1_w = main_nist_clock_nist_clock_timer0_reload_storage_full[15:8];
assign builder_nist_clock_csrbank13_reload0_w = main_nist_clock_nist_clock_timer0_reload_storage_full[7:0];
assign main_nist_clock_nist_clock_timer0_en_storage = main_nist_clock_nist_clock_timer0_en_storage_full;
assign builder_nist_clock_csrbank13_en0_w = main_nist_clock_nist_clock_timer0_en_storage_full;
assign builder_nist_clock_csrbank13_value7_w = main_nist_clock_nist_clock_timer0_value_status[63:56];
assign builder_nist_clock_csrbank13_value6_w = main_nist_clock_nist_clock_timer0_value_status[55:48];
assign builder_nist_clock_csrbank13_value5_w = main_nist_clock_nist_clock_timer0_value_status[47:40];
assign builder_nist_clock_csrbank13_value4_w = main_nist_clock_nist_clock_timer0_value_status[39:32];
assign builder_nist_clock_csrbank13_value3_w = main_nist_clock_nist_clock_timer0_value_status[31:24];
assign builder_nist_clock_csrbank13_value2_w = main_nist_clock_nist_clock_timer0_value_status[23:16];
assign builder_nist_clock_csrbank13_value1_w = main_nist_clock_nist_clock_timer0_value_status[15:8];
assign builder_nist_clock_csrbank13_value0_w = main_nist_clock_nist_clock_timer0_value_status[7:0];
assign main_nist_clock_nist_clock_timer0_eventmanager_storage = main_nist_clock_nist_clock_timer0_eventmanager_storage_full;
assign builder_nist_clock_csrbank13_ev_enable0_w = main_nist_clock_nist_clock_timer0_eventmanager_storage_full;
assign builder_nist_clock_csrbank14_sel = (builder_nist_clock_interface14_bank_bus_adr[13:9] == 4'd12);
assign builder_nist_clock_csrbank14_load7_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load7_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 1'd0));
assign builder_nist_clock_csrbank14_load6_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load6_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 1'd1));
assign builder_nist_clock_csrbank14_load5_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load5_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 2'd2));
assign builder_nist_clock_csrbank14_load4_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load4_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 2'd3));
assign builder_nist_clock_csrbank14_load3_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load3_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 3'd4));
assign builder_nist_clock_csrbank14_load2_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load2_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 3'd5));
assign builder_nist_clock_csrbank14_load1_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load1_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 3'd6));
assign builder_nist_clock_csrbank14_load0_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_load0_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 3'd7));
assign builder_nist_clock_csrbank14_reload7_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload7_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd8));
assign builder_nist_clock_csrbank14_reload6_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload6_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd9));
assign builder_nist_clock_csrbank14_reload5_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload5_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd10));
assign builder_nist_clock_csrbank14_reload4_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload4_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd11));
assign builder_nist_clock_csrbank14_reload3_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload3_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd12));
assign builder_nist_clock_csrbank14_reload2_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload2_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd13));
assign builder_nist_clock_csrbank14_reload1_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload1_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd14));
assign builder_nist_clock_csrbank14_reload0_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_reload0_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 4'd15));
assign builder_nist_clock_csrbank14_en0_r = builder_nist_clock_interface14_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank14_en0_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd16));
assign main_update_value_r = builder_nist_clock_interface14_bank_bus_dat_w[0];
assign main_update_value_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd17));
assign builder_nist_clock_csrbank14_value7_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value7_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd18));
assign builder_nist_clock_csrbank14_value6_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value6_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd19));
assign builder_nist_clock_csrbank14_value5_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value5_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd20));
assign builder_nist_clock_csrbank14_value4_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value4_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd21));
assign builder_nist_clock_csrbank14_value3_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value3_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd22));
assign builder_nist_clock_csrbank14_value2_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value2_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd23));
assign builder_nist_clock_csrbank14_value1_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value1_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd24));
assign builder_nist_clock_csrbank14_value0_r = builder_nist_clock_interface14_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank14_value0_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd25));
assign main_eventmanager_status_r = builder_nist_clock_interface14_bank_bus_dat_w[0];
assign main_eventmanager_status_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd26));
assign main_eventmanager_pending_r = builder_nist_clock_interface14_bank_bus_dat_w[0];
assign main_eventmanager_pending_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd27));
assign builder_nist_clock_csrbank14_ev_enable0_r = builder_nist_clock_interface14_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank14_ev_enable0_re = ((builder_nist_clock_csrbank14_sel & builder_nist_clock_interface14_bank_bus_we) & (builder_nist_clock_interface14_bank_bus_adr[4:0] == 5'd28));
assign main_load_storage = main_load_storage_full[63:0];
assign builder_nist_clock_csrbank14_load7_w = main_load_storage_full[63:56];
assign builder_nist_clock_csrbank14_load6_w = main_load_storage_full[55:48];
assign builder_nist_clock_csrbank14_load5_w = main_load_storage_full[47:40];
assign builder_nist_clock_csrbank14_load4_w = main_load_storage_full[39:32];
assign builder_nist_clock_csrbank14_load3_w = main_load_storage_full[31:24];
assign builder_nist_clock_csrbank14_load2_w = main_load_storage_full[23:16];
assign builder_nist_clock_csrbank14_load1_w = main_load_storage_full[15:8];
assign builder_nist_clock_csrbank14_load0_w = main_load_storage_full[7:0];
assign main_reload_storage = main_reload_storage_full[63:0];
assign builder_nist_clock_csrbank14_reload7_w = main_reload_storage_full[63:56];
assign builder_nist_clock_csrbank14_reload6_w = main_reload_storage_full[55:48];
assign builder_nist_clock_csrbank14_reload5_w = main_reload_storage_full[47:40];
assign builder_nist_clock_csrbank14_reload4_w = main_reload_storage_full[39:32];
assign builder_nist_clock_csrbank14_reload3_w = main_reload_storage_full[31:24];
assign builder_nist_clock_csrbank14_reload2_w = main_reload_storage_full[23:16];
assign builder_nist_clock_csrbank14_reload1_w = main_reload_storage_full[15:8];
assign builder_nist_clock_csrbank14_reload0_w = main_reload_storage_full[7:0];
assign main_en_storage = main_en_storage_full;
assign builder_nist_clock_csrbank14_en0_w = main_en_storage_full;
assign builder_nist_clock_csrbank14_value7_w = main_value_status[63:56];
assign builder_nist_clock_csrbank14_value6_w = main_value_status[55:48];
assign builder_nist_clock_csrbank14_value5_w = main_value_status[47:40];
assign builder_nist_clock_csrbank14_value4_w = main_value_status[39:32];
assign builder_nist_clock_csrbank14_value3_w = main_value_status[31:24];
assign builder_nist_clock_csrbank14_value2_w = main_value_status[23:16];
assign builder_nist_clock_csrbank14_value1_w = main_value_status[15:8];
assign builder_nist_clock_csrbank14_value0_w = main_value_status[7:0];
assign main_eventmanager_storage = main_eventmanager_storage_full;
assign builder_nist_clock_csrbank14_ev_enable0_w = main_eventmanager_storage_full;
assign builder_nist_clock_csrbank15_sel = (builder_nist_clock_interface15_bank_bus_adr[13:9] == 3'd4);
assign builder_nist_clock_csrbank15_enable_null0_r = builder_nist_clock_interface15_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank15_enable_null0_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 1'd0));
assign builder_nist_clock_csrbank15_enable_prog0_r = builder_nist_clock_interface15_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank15_enable_prog0_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 1'd1));
assign builder_nist_clock_csrbank15_prog_address3_r = builder_nist_clock_interface15_bank_bus_dat_w[5:0];
assign builder_nist_clock_csrbank15_prog_address3_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 2'd2));
assign builder_nist_clock_csrbank15_prog_address2_r = builder_nist_clock_interface15_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank15_prog_address2_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 2'd3));
assign builder_nist_clock_csrbank15_prog_address1_r = builder_nist_clock_interface15_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank15_prog_address1_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 3'd4));
assign builder_nist_clock_csrbank15_prog_address0_r = builder_nist_clock_interface15_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank15_prog_address0_re = ((builder_nist_clock_csrbank15_sel & builder_nist_clock_interface15_bank_bus_we) & (builder_nist_clock_interface15_bank_bus_adr[2:0] == 3'd5));
assign main_nist_clock_nist_clock_tmpu_enable_null_storage = main_nist_clock_nist_clock_tmpu_enable_null_storage_full;
assign builder_nist_clock_csrbank15_enable_null0_w = main_nist_clock_nist_clock_tmpu_enable_null_storage_full;
assign main_nist_clock_nist_clock_tmpu_enable_prog_storage = main_nist_clock_nist_clock_tmpu_enable_prog_storage_full;
assign builder_nist_clock_csrbank15_enable_prog0_w = main_nist_clock_nist_clock_tmpu_enable_prog_storage_full;
assign main_nist_clock_nist_clock_tmpu_prog_address_storage = main_nist_clock_nist_clock_tmpu_prog_address_storage_full[29:12];
assign builder_nist_clock_csrbank15_prog_address3_w = main_nist_clock_nist_clock_tmpu_prog_address_storage_full[29:24];
assign builder_nist_clock_csrbank15_prog_address2_w = main_nist_clock_nist_clock_tmpu_prog_address_storage_full[23:16];
assign builder_nist_clock_csrbank15_prog_address1_w = {main_nist_clock_nist_clock_tmpu_prog_address_storage_full[15:12], {4{1'd0}}};
assign builder_nist_clock_csrbank15_prog_address0_w = 1'd0;
assign builder_nist_clock_csrbank16_sel = (builder_nist_clock_interface16_bank_bus_adr[13:9] == 1'd1);
assign main_nist_clock_nist_clock_uart_rxtx_r = builder_nist_clock_interface16_bank_bus_dat_w[7:0];
assign main_nist_clock_nist_clock_uart_rxtx_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 1'd0));
assign builder_nist_clock_csrbank16_txfull_r = builder_nist_clock_interface16_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank16_txfull_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 1'd1));
assign builder_nist_clock_csrbank16_rxempty_r = builder_nist_clock_interface16_bank_bus_dat_w[0];
assign builder_nist_clock_csrbank16_rxempty_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 2'd2));
assign main_nist_clock_nist_clock_uart_status_r = builder_nist_clock_interface16_bank_bus_dat_w[1:0];
assign main_nist_clock_nist_clock_uart_status_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 2'd3));
assign main_nist_clock_nist_clock_uart_pending_r = builder_nist_clock_interface16_bank_bus_dat_w[1:0];
assign main_nist_clock_nist_clock_uart_pending_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 3'd4));
assign builder_nist_clock_csrbank16_ev_enable0_r = builder_nist_clock_interface16_bank_bus_dat_w[1:0];
assign builder_nist_clock_csrbank16_ev_enable0_re = ((builder_nist_clock_csrbank16_sel & builder_nist_clock_interface16_bank_bus_we) & (builder_nist_clock_interface16_bank_bus_adr[2:0] == 3'd5));
assign builder_nist_clock_csrbank16_txfull_w = main_nist_clock_nist_clock_uart_txfull_status;
assign builder_nist_clock_csrbank16_rxempty_w = main_nist_clock_nist_clock_uart_rxempty_status;
assign main_nist_clock_nist_clock_uart_storage = main_nist_clock_nist_clock_uart_storage_full[1:0];
assign builder_nist_clock_csrbank16_ev_enable0_w = main_nist_clock_nist_clock_uart_storage_full[1:0];
assign builder_nist_clock_csrbank17_sel = (builder_nist_clock_interface17_bank_bus_adr[13:9] == 1'd0);
assign builder_nist_clock_csrbank17_tuning_word3_r = builder_nist_clock_interface17_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank17_tuning_word3_re = ((builder_nist_clock_csrbank17_sel & builder_nist_clock_interface17_bank_bus_we) & (builder_nist_clock_interface17_bank_bus_adr[1:0] == 1'd0));
assign builder_nist_clock_csrbank17_tuning_word2_r = builder_nist_clock_interface17_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank17_tuning_word2_re = ((builder_nist_clock_csrbank17_sel & builder_nist_clock_interface17_bank_bus_we) & (builder_nist_clock_interface17_bank_bus_adr[1:0] == 1'd1));
assign builder_nist_clock_csrbank17_tuning_word1_r = builder_nist_clock_interface17_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank17_tuning_word1_re = ((builder_nist_clock_csrbank17_sel & builder_nist_clock_interface17_bank_bus_we) & (builder_nist_clock_interface17_bank_bus_adr[1:0] == 2'd2));
assign builder_nist_clock_csrbank17_tuning_word0_r = builder_nist_clock_interface17_bank_bus_dat_w[7:0];
assign builder_nist_clock_csrbank17_tuning_word0_re = ((builder_nist_clock_csrbank17_sel & builder_nist_clock_interface17_bank_bus_we) & (builder_nist_clock_interface17_bank_bus_adr[1:0] == 2'd3));
assign main_nist_clock_nist_clock_uart_phy_storage = main_nist_clock_nist_clock_uart_phy_storage_full[31:0];
assign builder_nist_clock_csrbank17_tuning_word3_w = main_nist_clock_nist_clock_uart_phy_storage_full[31:24];
assign builder_nist_clock_csrbank17_tuning_word2_w = main_nist_clock_nist_clock_uart_phy_storage_full[23:16];
assign builder_nist_clock_csrbank17_tuning_word1_w = main_nist_clock_nist_clock_uart_phy_storage_full[15:8];
assign builder_nist_clock_csrbank17_tuning_word0_w = main_nist_clock_nist_clock_uart_phy_storage_full[7:0];
assign builder_nist_clock_interface0_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface1_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface2_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface3_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface4_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface5_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface6_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface7_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface8_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface9_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface10_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface11_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface12_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface13_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface14_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface15_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface16_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface17_bank_bus_adr = main_nist_clock_nist_clock_interface_adr;
assign builder_nist_clock_interface0_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface1_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface2_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface3_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface4_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface5_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface6_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface7_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface8_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface9_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface10_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface11_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface12_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface13_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface14_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface15_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface16_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface17_bank_bus_we = main_nist_clock_nist_clock_interface_we;
assign builder_nist_clock_interface0_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface1_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface2_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface3_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface4_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface5_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface6_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface7_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface8_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface9_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface10_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface11_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface12_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface13_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface14_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface15_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface16_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign builder_nist_clock_interface17_bank_bus_dat_w = main_nist_clock_nist_clock_interface_dat_w;
assign main_nist_clock_nist_clock_interface_dat_r = (((((((((((((((((builder_nist_clock_interface0_bank_bus_dat_r | builder_nist_clock_interface1_bank_bus_dat_r) | builder_nist_clock_interface2_bank_bus_dat_r) | builder_nist_clock_interface3_bank_bus_dat_r) | builder_nist_clock_interface4_bank_bus_dat_r) | builder_nist_clock_interface5_bank_bus_dat_r) | builder_nist_clock_interface6_bank_bus_dat_r) | builder_nist_clock_interface7_bank_bus_dat_r) | builder_nist_clock_interface8_bank_bus_dat_r) | builder_nist_clock_interface9_bank_bus_dat_r) | builder_nist_clock_interface10_bank_bus_dat_r) | builder_nist_clock_interface11_bank_bus_dat_r) | builder_nist_clock_interface12_bank_bus_dat_r) | builder_nist_clock_interface13_bank_bus_dat_r) | builder_nist_clock_interface14_bank_bus_dat_r) | builder_nist_clock_interface15_bank_bus_dat_r) | builder_nist_clock_interface16_bank_bus_dat_r) | builder_nist_clock_interface17_bank_bus_dat_r);

// synthesis translate_off
reg dummy_d_174;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed0 <= 30'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed0 <= main_kernel_cpu_ibus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed0 <= main_kernel_cpu_dbus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_174 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_175;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed1 <= 32'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed1 <= main_kernel_cpu_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed1 <= main_kernel_cpu_dbus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_175 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_176;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed2 <= 4'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed2 <= main_kernel_cpu_ibus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed2 <= main_kernel_cpu_dbus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_176 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_177;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed3 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed3 <= main_kernel_cpu_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed3 <= main_kernel_cpu_dbus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_177 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_178;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed4 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed4 <= main_kernel_cpu_ibus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed4 <= main_kernel_cpu_dbus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_178 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_179;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed5 <= 1'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed5 <= main_kernel_cpu_ibus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed5 <= main_kernel_cpu_dbus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_179 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_180;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed6 <= 3'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed6 <= main_kernel_cpu_ibus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed6 <= main_kernel_cpu_dbus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_180 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_181;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed7 <= 2'd0;
	case (builder_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed7 <= main_kernel_cpu_ibus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed7 <= main_kernel_cpu_dbus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_181 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_182;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed8 <= 1'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record0_writable;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record1_writable;
		end
		2'd2: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record2_writable;
		end
		2'd3: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record3_writable;
		end
		3'd4: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record4_writable;
		end
		3'd5: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record5_writable;
		end
		3'd6: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record6_writable;
		end
		default: begin
			builder_comb_rhs_array_muxed8 <= main_rtio_core_outputs_lanedistributor_record7_writable;
		end
	endcase
// synthesis translate_off
	dummy_d_182 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_183;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed9 <= 2'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		2'd2: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		2'd3: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow0, (main_rtio_core_inputs_asyncfifo0_asyncfifo0_readable & (~main_rtio_core_inputs_overflow0))};
		end
		3'd4: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd5: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd6: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		3'd7: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow1, (main_rtio_core_inputs_asyncfifo1_asyncfifo1_readable & (~main_rtio_core_inputs_overflow1))};
		end
		4'd8: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd9: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd10: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd11: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow2, (main_rtio_core_inputs_asyncfifo2_asyncfifo2_readable & (~main_rtio_core_inputs_overflow2))};
		end
		4'd12: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd13: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd14: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		4'd15: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow3, (main_rtio_core_inputs_asyncfifo3_asyncfifo3_readable & (~main_rtio_core_inputs_overflow3))};
		end
		5'd16: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow4, (main_rtio_core_inputs_asyncfifo4_asyncfifo4_readable & (~main_rtio_core_inputs_overflow4))};
		end
		5'd17: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow5, (main_rtio_core_inputs_asyncfifo5_asyncfifo5_readable & (~main_rtio_core_inputs_overflow5))};
		end
		5'd18: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow6, (main_rtio_core_inputs_asyncfifo6_asyncfifo6_readable & (~main_rtio_core_inputs_overflow6))};
		end
		5'd19: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd20: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd21: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		5'd22: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow7, (main_rtio_core_inputs_asyncfifo7_asyncfifo7_readable & (~main_rtio_core_inputs_overflow7))};
		end
		5'd23: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow8, (main_rtio_core_inputs_asyncfifo8_asyncfifo8_readable & (~main_rtio_core_inputs_overflow8))};
		end
		5'd24: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow9, (main_rtio_core_inputs_asyncfifo9_asyncfifo9_readable & (~main_rtio_core_inputs_overflow9))};
		end
		5'd25: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow10, (main_rtio_core_inputs_asyncfifo10_asyncfifo10_readable & (~main_rtio_core_inputs_overflow10))};
		end
		5'd26: begin
			builder_comb_rhs_array_muxed9 <= {main_rtio_core_inputs_overflow11, (main_rtio_core_inputs_asyncfifo11_asyncfifo11_readable & (~main_rtio_core_inputs_overflow11))};
		end
		5'd27: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_183 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_184;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed10 <= 2'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed10 <= main_rtio_cri_cmd;
		end
		default: begin
			builder_comb_rhs_array_muxed10 <= main_dma_cri_master_cri_cmd;
		end
	endcase
// synthesis translate_off
	dummy_d_184 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_185;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed11 <= 24'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed11 <= main_rtio_cri_chan_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed11 <= main_dma_cri_master_cri_chan_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_185 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_186;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed12 <= 64'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed12 <= main_rtio_cri_o_timestamp;
		end
		default: begin
			builder_comb_rhs_array_muxed12 <= main_dma_cri_master_cri_o_timestamp;
		end
	endcase
// synthesis translate_off
	dummy_d_186 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_187;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed13 <= 512'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed13 <= main_rtio_cri_o_data;
		end
		default: begin
			builder_comb_rhs_array_muxed13 <= main_dma_cri_master_cri_o_data;
		end
	endcase
// synthesis translate_off
	dummy_d_187 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_188;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed14 <= 8'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed14 <= main_rtio_cri_o_address;
		end
		default: begin
			builder_comb_rhs_array_muxed14 <= main_dma_cri_master_cri_o_address;
		end
	endcase
// synthesis translate_off
	dummy_d_188 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_189;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed15 <= 64'd0;
	case (main_cri_con_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed15 <= main_rtio_cri_i_timeout;
		end
		default: begin
			builder_comb_rhs_array_muxed15 <= main_dma_cri_master_cri_i_timeout;
		end
	endcase
// synthesis translate_off
	dummy_d_189 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_190;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed17 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed17 <= main_inj_o_sys0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed17 <= main_inj_o_sys1;
		end
		default: begin
			builder_comb_rhs_array_muxed17 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_190 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_191;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed18 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed18 <= main_inj_o_sys2;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed18 <= main_inj_o_sys3;
		end
		default: begin
			builder_comb_rhs_array_muxed18 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_191 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_192;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed19 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed19 <= main_inj_o_sys4;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed19 <= main_inj_o_sys5;
		end
		default: begin
			builder_comb_rhs_array_muxed19 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_192 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_193;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed20 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys6;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys7;
		end
		default: begin
			builder_comb_rhs_array_muxed20 <= main_inj_o_sys8;
		end
	endcase
// synthesis translate_off
	dummy_d_193 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_194;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed21 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed21 <= main_inj_o_sys9;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed21 <= main_inj_o_sys10;
		end
		default: begin
			builder_comb_rhs_array_muxed21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_194 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_195;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed22 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed22 <= main_inj_o_sys11;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed22 <= main_inj_o_sys12;
		end
		default: begin
			builder_comb_rhs_array_muxed22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_195 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_196;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed23 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed23 <= main_inj_o_sys13;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed23 <= main_inj_o_sys14;
		end
		default: begin
			builder_comb_rhs_array_muxed23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_196 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_197;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed24 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys15;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys16;
		end
		default: begin
			builder_comb_rhs_array_muxed24 <= main_inj_o_sys17;
		end
	endcase
// synthesis translate_off
	dummy_d_197 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_198;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed25 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed25 <= main_inj_o_sys18;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed25 <= main_inj_o_sys19;
		end
		default: begin
			builder_comb_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_198 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_199;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed26 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed26 <= main_inj_o_sys20;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed26 <= main_inj_o_sys21;
		end
		default: begin
			builder_comb_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_199 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_200;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed27 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed27 <= main_inj_o_sys22;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed27 <= main_inj_o_sys23;
		end
		default: begin
			builder_comb_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_200 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_201;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed28 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed28 <= main_inj_o_sys24;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed28 <= main_inj_o_sys25;
		end
		default: begin
			builder_comb_rhs_array_muxed28 <= main_inj_o_sys26;
		end
	endcase
// synthesis translate_off
	dummy_d_201 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_202;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed29 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed29 <= main_inj_o_sys27;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed29 <= main_inj_o_sys28;
		end
		default: begin
			builder_comb_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_202 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_203;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed30 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed30 <= main_inj_o_sys29;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed30 <= main_inj_o_sys30;
		end
		default: begin
			builder_comb_rhs_array_muxed30 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_203 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_204;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed31 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed31 <= main_inj_o_sys31;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed31 <= main_inj_o_sys32;
		end
		default: begin
			builder_comb_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_204 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_205;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed32 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed32 <= main_inj_o_sys33;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed32 <= main_inj_o_sys34;
		end
		default: begin
			builder_comb_rhs_array_muxed32 <= main_inj_o_sys35;
		end
	endcase
// synthesis translate_off
	dummy_d_205 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_206;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed33 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed33 <= main_inj_o_sys36;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed33 <= main_inj_o_sys37;
		end
		default: begin
			builder_comb_rhs_array_muxed33 <= main_inj_o_sys38;
		end
	endcase
// synthesis translate_off
	dummy_d_206 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_207;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed34 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed34 <= main_inj_o_sys39;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed34 <= main_inj_o_sys40;
		end
		default: begin
			builder_comb_rhs_array_muxed34 <= main_inj_o_sys41;
		end
	endcase
// synthesis translate_off
	dummy_d_207 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_208;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed35 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed35 <= main_inj_o_sys42;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed35 <= main_inj_o_sys43;
		end
		default: begin
			builder_comb_rhs_array_muxed35 <= main_inj_o_sys44;
		end
	endcase
// synthesis translate_off
	dummy_d_208 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_209;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed36 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed36 <= main_inj_o_sys45;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed36 <= main_inj_o_sys46;
		end
		default: begin
			builder_comb_rhs_array_muxed36 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_209 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_210;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed37 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed37 <= main_inj_o_sys47;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed37 <= main_inj_o_sys48;
		end
		default: begin
			builder_comb_rhs_array_muxed37 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_210 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_211;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed38 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed38 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed38 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed38 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_211 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_212;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed39 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed39 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_212 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_213;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed40 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed40 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed40 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed40 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_213 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_214;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed41 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed41 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed41 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed41 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_214 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_215;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed42 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed42 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed42 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed42 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_215 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_216;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed43 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed43 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed43 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed43 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_216 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_217;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed44 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed44 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed44 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed44 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_217 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_218;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed45 <= 1'd0;
	case (main_inj_override_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
		default: begin
			builder_comb_rhs_array_muxed45 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_218 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_219;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed16 <= 1'd0;
	case (main_inj_chan_sel_storage)
		1'd0: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed17;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed18;
		end
		2'd2: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed19;
		end
		2'd3: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed20;
		end
		3'd4: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed21;
		end
		3'd5: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed22;
		end
		3'd6: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed23;
		end
		3'd7: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed24;
		end
		4'd8: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed25;
		end
		4'd9: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed26;
		end
		4'd10: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed27;
		end
		4'd11: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed28;
		end
		4'd12: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed29;
		end
		4'd13: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed30;
		end
		4'd14: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed31;
		end
		4'd15: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed32;
		end
		5'd16: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed33;
		end
		5'd17: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed34;
		end
		5'd18: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed35;
		end
		5'd19: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed36;
		end
		5'd20: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed37;
		end
		5'd21: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed38;
		end
		5'd22: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed39;
		end
		5'd23: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed40;
		end
		5'd24: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed41;
		end
		5'd25: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed42;
		end
		5'd26: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed43;
		end
		5'd27: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed44;
		end
		default: begin
			builder_comb_rhs_array_muxed16 <= builder_comb_rhs_array_muxed45;
		end
	endcase
// synthesis translate_off
	dummy_d_219 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_220;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed46 <= 30'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed46 <= main_nist_clock_nist_clock_wb_sdram_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed46 <= main_kernel_cpu_wb_sdram_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_220 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_221;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed47 <= 32'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed47 <= main_nist_clock_nist_clock_wb_sdram_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed47 <= main_kernel_cpu_wb_sdram_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_221 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_222;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed48 <= 4'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed48 <= main_nist_clock_nist_clock_wb_sdram_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed48 <= main_kernel_cpu_wb_sdram_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_222 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_223;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed49 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed49 <= main_nist_clock_nist_clock_wb_sdram_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed49 <= main_kernel_cpu_wb_sdram_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_223 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_224;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed50 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed50 <= main_nist_clock_nist_clock_wb_sdram_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed50 <= main_kernel_cpu_wb_sdram_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_224 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_225;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed51 <= 1'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed51 <= main_nist_clock_nist_clock_wb_sdram_we;
		end
		default: begin
			builder_comb_rhs_array_muxed51 <= main_kernel_cpu_wb_sdram_we;
		end
	endcase
// synthesis translate_off
	dummy_d_225 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_226;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed52 <= 3'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed52 <= main_nist_clock_nist_clock_wb_sdram_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed52 <= main_kernel_cpu_wb_sdram_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_226 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_227;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed53 <= 2'd0;
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed53 <= main_nist_clock_nist_clock_wb_sdram_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed53 <= main_kernel_cpu_wb_sdram_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_227 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_228;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed54 <= 30'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed54 <= main_nist_clock_nist_clock_bridge_if_bus_adr;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed54 <= main_interface0_bus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed54 <= main_interface1_bus_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_228 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_229;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed55 <= 512'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed55 <= main_nist_clock_nist_clock_bridge_if_bus_dat_w;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed55 <= main_interface0_bus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed55 <= main_interface1_bus_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_229 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_230;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed56 <= 64'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed56 <= main_nist_clock_nist_clock_bridge_if_bus_sel;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed56 <= main_interface0_bus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed56 <= main_interface1_bus_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_230 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_231;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed57 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed57 <= main_nist_clock_nist_clock_bridge_if_bus_cyc;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed57 <= main_interface0_bus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed57 <= main_interface1_bus_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_231 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_232;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed58 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed58 <= main_nist_clock_nist_clock_bridge_if_bus_stb;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed58 <= main_interface0_bus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed58 <= main_interface1_bus_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_232 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_233;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed59 <= 1'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed59 <= main_nist_clock_nist_clock_bridge_if_bus_we;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed59 <= main_interface0_bus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed59 <= main_interface1_bus_we;
		end
	endcase
// synthesis translate_off
	dummy_d_233 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_234;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed60 <= 3'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed60 <= main_nist_clock_nist_clock_bridge_if_bus_cti;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed60 <= main_interface0_bus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed60 <= main_interface1_bus_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_234 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_235;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed61 <= 2'd0;
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed61 <= main_nist_clock_nist_clock_bridge_if_bus_bte;
		end
		1'd1: begin
			builder_comb_rhs_array_muxed61 <= main_interface0_bus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed61 <= main_interface1_bus_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_235 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_236;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed62 <= 30'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed62 <= main_nist_clock_nist_clock_ibus_adr;
		end
		default: begin
			builder_comb_rhs_array_muxed62 <= main_nist_clock_nist_clock_tmpu_adr;
		end
	endcase
// synthesis translate_off
	dummy_d_236 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_237;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed63 <= 32'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed63 <= main_nist_clock_nist_clock_ibus_dat_w;
		end
		default: begin
			builder_comb_rhs_array_muxed63 <= main_nist_clock_nist_clock_tmpu_dat_w;
		end
	endcase
// synthesis translate_off
	dummy_d_237 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_238;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed64 <= 4'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed64 <= main_nist_clock_nist_clock_ibus_sel;
		end
		default: begin
			builder_comb_rhs_array_muxed64 <= main_nist_clock_nist_clock_tmpu_sel;
		end
	endcase
// synthesis translate_off
	dummy_d_238 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_239;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed65 <= 1'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed65 <= main_nist_clock_nist_clock_ibus_cyc;
		end
		default: begin
			builder_comb_rhs_array_muxed65 <= main_nist_clock_nist_clock_tmpu_cyc;
		end
	endcase
// synthesis translate_off
	dummy_d_239 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_240;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed66 <= 1'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed66 <= main_nist_clock_nist_clock_ibus_stb;
		end
		default: begin
			builder_comb_rhs_array_muxed66 <= main_nist_clock_nist_clock_tmpu_stb;
		end
	endcase
// synthesis translate_off
	dummy_d_240 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_241;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed67 <= 1'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed67 <= main_nist_clock_nist_clock_ibus_we;
		end
		default: begin
			builder_comb_rhs_array_muxed67 <= main_nist_clock_nist_clock_tmpu_we;
		end
	endcase
// synthesis translate_off
	dummy_d_241 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_242;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed68 <= 3'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed68 <= main_nist_clock_nist_clock_ibus_cti;
		end
		default: begin
			builder_comb_rhs_array_muxed68 <= main_nist_clock_nist_clock_tmpu_cti;
		end
	endcase
// synthesis translate_off
	dummy_d_242 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_243;
// synthesis translate_on
always @(*) begin
	builder_comb_rhs_array_muxed69 <= 2'd0;
	case (builder_nist_clock_grant)
		1'd0: begin
			builder_comb_rhs_array_muxed69 <= main_nist_clock_nist_clock_ibus_bte;
		end
		default: begin
			builder_comb_rhs_array_muxed69 <= main_nist_clock_nist_clock_tmpu_bte;
		end
	endcase
// synthesis translate_off
	dummy_d_243 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_244;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed0 <= 1'd0;
	case (main_rtio_core_outputs_channel_r0)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed0 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed0 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed0 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed0 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed0 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed0 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_244 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_245;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed1 <= 1'd0;
	case (main_rtio_core_outputs_channel_r1)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed1 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed1 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed1 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed1 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed1 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed1 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_245 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_246;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed2 <= 1'd0;
	case (main_rtio_core_outputs_channel_r2)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed2 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed2 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed2 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed2 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed2 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed2 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_246 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_247;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed3 <= 1'd0;
	case (main_rtio_core_outputs_channel_r3)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed3 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed3 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed3 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed3 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed3 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed3 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_247 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_248;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed4 <= 1'd0;
	case (main_rtio_core_outputs_channel_r4)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed4 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed4 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed4 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed4 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed4 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed4 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_248 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_249;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed5 <= 1'd0;
	case (main_rtio_core_outputs_channel_r5)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed5 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed5 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed5 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed5 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed5 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed5 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_249 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_250;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed6 <= 1'd0;
	case (main_rtio_core_outputs_channel_r6)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed6 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed6 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed6 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed6 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed6 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed6 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_250 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_251;
// synthesis translate_on
always @(*) begin
	builder_sync_basiclowerer_array_muxed7 <= 1'd0;
	case (main_rtio_core_outputs_channel_r7)
		1'd0: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x0_busy;
		end
		1'd1: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x1_busy;
		end
		2'd2: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x2_busy;
		end
		2'd3: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x0_inout_8x0_ointerface0_busy;
		end
		3'd4: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x3_busy;
		end
		3'd5: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x4_busy;
		end
		3'd6: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x5_busy;
		end
		3'd7: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x1_inout_8x1_ointerface1_busy;
		end
		4'd8: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x6_busy;
		end
		4'd9: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x7_busy;
		end
		4'd10: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x8_busy;
		end
		4'd11: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x2_inout_8x2_ointerface2_busy;
		end
		4'd12: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x9_busy;
		end
		4'd13: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x10_busy;
		end
		4'd14: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output_8x11_busy;
		end
		4'd15: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x3_inout_8x3_ointerface3_busy;
		end
		5'd16: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x4_inout_8x4_ointerface4_busy;
		end
		5'd17: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x5_inout_8x5_ointerface5_busy;
		end
		5'd18: begin
			builder_sync_basiclowerer_array_muxed7 <= main_inout_8x6_inout_8x6_ointerface6_busy;
		end
		5'd19: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output0_busy;
		end
		5'd20: begin
			builder_sync_basiclowerer_array_muxed7 <= main_output1_busy;
		end
		5'd21: begin
			builder_sync_basiclowerer_array_muxed7 <= main_clockgen_busy;
		end
		5'd22: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster0_ointerface0_busy;
		end
		5'd23: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster1_ointerface1_busy;
		end
		5'd24: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster2_ointerface2_busy;
		end
		5'd25: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster3_ointerface3_busy;
		end
		5'd26: begin
			builder_sync_basiclowerer_array_muxed7 <= main_spimaster4_ointerface4_busy;
		end
		5'd27: begin
			builder_sync_basiclowerer_array_muxed7 <= main_ad9914_busy;
		end
		default: begin
			builder_sync_basiclowerer_array_muxed7 <= main_busy;
		end
	endcase
// synthesis translate_off
	dummy_d_251 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_252;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed0 <= 8'd0;
	case (main_output_8x0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed0 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed0 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed0 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed0 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed0 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed0 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed0 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed0 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_252 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_253;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed0 <= 7'd0;
	case (main_output_8x0_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed0 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed0 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed0 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed0 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed0 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed0 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed0 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_253 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_254;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed1 <= 8'd0;
	case (main_output_8x1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed1 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed1 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed1 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed1 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed1 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed1 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed1 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed1 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_254 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_255;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed1 <= 7'd0;
	case (main_output_8x1_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed1 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed1 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed1 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed1 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed1 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed1 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed1 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed1 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_255 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_256;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed2 <= 8'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed2 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed2 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed2 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed2 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed2 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed2 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed2 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed2 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_256 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_257;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed2 <= 7'd0;
	case (main_output_8x2_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed2 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed2 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed2 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed2 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed2 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed2 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed2 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed2 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_257 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_258;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed3 <= 8'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed3 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed3 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed3 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed3 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed3 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed3 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed3 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed3 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_258 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_259;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed3 <= 7'd0;
	case (main_inout_8x0_inout_8x0_ointerface0_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed3 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed3 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed3 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed3 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed3 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed3 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed3 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed3 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_259 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_260;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed4 <= 8'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed4 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed4 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed4 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed4 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed4 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed4 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed4 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed4 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_260 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_261;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed4 <= 7'd0;
	case (main_output_8x3_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed4 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed4 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed4 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed4 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed4 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed4 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed4 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed4 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_261 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_262;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed5 <= 8'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed5 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed5 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed5 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed5 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed5 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed5 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed5 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed5 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_262 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_263;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed5 <= 7'd0;
	case (main_output_8x4_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed5 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed5 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed5 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed5 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed5 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed5 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed5 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed5 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_263 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_264;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed6 <= 8'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed6 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed6 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed6 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed6 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed6 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed6 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed6 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed6 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_264 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_265;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed6 <= 7'd0;
	case (main_output_8x5_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed6 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed6 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed6 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed6 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed6 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed6 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed6 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_265 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_266;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed7 <= 8'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed7 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed7 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed7 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed7 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed7 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed7 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed7 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed7 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_266 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_267;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed7 <= 7'd0;
	case (main_inout_8x1_inout_8x1_ointerface1_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed7 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed7 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed7 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed7 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed7 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed7 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed7 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed7 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_267 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_268;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed8 <= 8'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed8 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed8 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed8 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed8 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed8 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed8 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed8 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed8 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_268 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_269;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed8 <= 7'd0;
	case (main_output_8x6_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed8 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed8 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed8 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed8 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed8 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed8 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed8 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed8 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_269 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_270;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed9 <= 8'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed9 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed9 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed9 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed9 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed9 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed9 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed9 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed9 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_270 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_271;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed9 <= 7'd0;
	case (main_output_8x7_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed9 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed9 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed9 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed9 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed9 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed9 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed9 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed9 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_271 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_272;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed10 <= 8'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed10 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed10 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed10 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed10 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed10 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed10 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed10 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed10 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_272 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_273;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed10 <= 7'd0;
	case (main_output_8x8_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed10 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed10 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed10 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed10 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed10 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed10 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed10 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed10 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_273 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_274;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed11 <= 8'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed11 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed11 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed11 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed11 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed11 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed11 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed11 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed11 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_274 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_275;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed11 <= 7'd0;
	case (main_inout_8x2_inout_8x2_ointerface2_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed11 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed11 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed11 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed11 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed11 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed11 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed11 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed11 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_275 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_276;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed12 <= 8'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed12 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed12 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed12 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed12 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed12 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed12 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed12 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed12 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_276 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_277;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed12 <= 7'd0;
	case (main_output_8x9_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed12 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed12 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed12 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed12 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed12 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed12 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed12 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_277 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_278;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed13 <= 8'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed13 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed13 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed13 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed13 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed13 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed13 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed13 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed13 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_278 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_279;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed13 <= 7'd0;
	case (main_output_8x10_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed13 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed13 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed13 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed13 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed13 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed13 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed13 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_279 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_280;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed14 <= 8'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed14 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed14 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed14 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed14 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed14 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed14 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed14 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed14 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_280 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_281;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed14 <= 7'd0;
	case (main_output_8x11_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed14 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed14 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed14 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed14 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed14 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed14 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed14 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed14 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_281 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_282;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed15 <= 8'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed15 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed15 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed15 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed15 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed15 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed15 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed15 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed15 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_282 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_283;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed15 <= 7'd0;
	case (main_inout_8x3_inout_8x3_ointerface3_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed15 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed15 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed15 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed15 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed15 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed15 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed15 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed15 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_283 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_284;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed16 <= 8'd0;
	case (main_inout_8x4_inout_8x4_ointerface4_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed16 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed16 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed16 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed16 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed16 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed16 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed16 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed16 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_284 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_285;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed16 <= 7'd0;
	case (main_inout_8x4_inout_8x4_ointerface4_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed16 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed16 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed16 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed16 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed16 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed16 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed16 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed16 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_285 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_286;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed17 <= 8'd0;
	case (main_inout_8x5_inout_8x5_ointerface5_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed17 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed17 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed17 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed17 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed17 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed17 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed17 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed17 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_286 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_287;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed17 <= 7'd0;
	case (main_inout_8x5_inout_8x5_ointerface5_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed17 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed17 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed17 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed17 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed17 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed17 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed17 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed17 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_287 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_288;
// synthesis translate_on
always @(*) begin
	builder_sync_f_t_array_muxed18 <= 8'd0;
	case (main_inout_8x6_inout_8x6_ointerface6_fine_ts)
		1'd0: begin
			builder_sync_f_t_array_muxed18 <= 8'd255;
		end
		1'd1: begin
			builder_sync_f_t_array_muxed18 <= 8'd254;
		end
		2'd2: begin
			builder_sync_f_t_array_muxed18 <= 8'd252;
		end
		2'd3: begin
			builder_sync_f_t_array_muxed18 <= 8'd248;
		end
		3'd4: begin
			builder_sync_f_t_array_muxed18 <= 8'd240;
		end
		3'd5: begin
			builder_sync_f_t_array_muxed18 <= 8'd224;
		end
		3'd6: begin
			builder_sync_f_t_array_muxed18 <= 8'd192;
		end
		default: begin
			builder_sync_f_t_array_muxed18 <= 8'd128;
		end
	endcase
// synthesis translate_off
	dummy_d_288 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_289;
// synthesis translate_on
always @(*) begin
	builder_sync_f_f_array_muxed18 <= 7'd0;
	case (main_inout_8x6_inout_8x6_ointerface6_fine_ts)
		1'd0: begin
			builder_sync_f_f_array_muxed18 <= 1'd0;
		end
		1'd1: begin
			builder_sync_f_f_array_muxed18 <= 1'd1;
		end
		2'd2: begin
			builder_sync_f_f_array_muxed18 <= 2'd3;
		end
		2'd3: begin
			builder_sync_f_f_array_muxed18 <= 3'd7;
		end
		3'd4: begin
			builder_sync_f_f_array_muxed18 <= 4'd15;
		end
		3'd5: begin
			builder_sync_f_f_array_muxed18 <= 5'd31;
		end
		3'd6: begin
			builder_sync_f_f_array_muxed18 <= 6'd63;
		end
		default: begin
			builder_sync_f_f_array_muxed18 <= 7'd127;
		end
	endcase
// synthesis translate_off
	dummy_d_289 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_290;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed0 <= 61'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane)
		1'd0: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			builder_sync_rhs_array_muxed0 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_290 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_291;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed1 <= 61'd0;
	case (main_rtio_core_outputs_lanedistributor_current_lane_plus_one)
		1'd0: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1;
		end
		2'd2: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2;
		end
		2'd3: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3;
		end
		3'd4: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4;
		end
		3'd5: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5;
		end
		3'd6: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6;
		end
		default: begin
			builder_sync_rhs_array_muxed1 <= main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7;
		end
	endcase
// synthesis translate_off
	dummy_d_291 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_292;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed0 <= 32'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record0_fifo_out_data;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record1_fifo_out_data;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record2_fifo_out_data;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record3_fifo_out_data;
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record4_fifo_out_data;
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record5_fifo_out_data;
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record6_fifo_out_data;
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record7_fifo_out_data;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record8_fifo_out_data;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record9_fifo_out_data;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record10_fifo_out_data;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed0 <= main_rtio_core_inputs_record11_fifo_out_data;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed0 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_292 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_293;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed1 <= 65'd0;
	case (main_rtio_core_cri_chan_sel[15:0])
		1'd0: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record0_fifo_out_timestamp <<< 1'd0);
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record1_fifo_out_timestamp <<< 1'd0);
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record2_fifo_out_timestamp <<< 1'd0);
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record3_fifo_out_timestamp <<< 1'd0);
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record4_fifo_out_timestamp <<< 1'd0);
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record5_fifo_out_timestamp <<< 1'd0);
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed1 <= (main_rtio_core_inputs_record6_fifo_out_timestamp <<< 1'd0);
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed1 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_293 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_294;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed2 <= 32'd0;
	case (main_mailbox_i1_adr[1:0])
		1'd0: begin
			builder_sync_rhs_array_muxed2 <= main_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed2 <= main_mailbox1;
		end
		default: begin
			builder_sync_rhs_array_muxed2 <= main_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_294 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_295;
// synthesis translate_on
always @(*) begin
	builder_sync_rhs_array_muxed3 <= 32'd0;
	case (main_mailbox_i2_adr[1:0])
		1'd0: begin
			builder_sync_rhs_array_muxed3 <= main_mailbox0;
		end
		1'd1: begin
			builder_sync_rhs_array_muxed3 <= main_mailbox1;
		end
		default: begin
			builder_sync_rhs_array_muxed3 <= main_mailbox2;
		end
	endcase
// synthesis translate_off
	dummy_d_295 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_296;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed3 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed3 <= main_mon_bussynchronizer0_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed3 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_296 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_297;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed4 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed4 <= main_mon_bussynchronizer1_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed4 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_297 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_298;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed5 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed5 <= main_mon_bussynchronizer2_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed5 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_298 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_299;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed6 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed6 <= main_mon_bussynchronizer3_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed6 <= main_mon_bussynchronizer4_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed6 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_299 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_300;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed7 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed7 <= main_mon_bussynchronizer5_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed7 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_300 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_301;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed8 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed8 <= main_mon_bussynchronizer6_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed8 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_301 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_302;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed9 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed9 <= main_mon_bussynchronizer7_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed9 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_302 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_303;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed10 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed10 <= main_mon_bussynchronizer8_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed10 <= main_mon_bussynchronizer9_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed10 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_303 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_304;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed11 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed11 <= main_mon_bussynchronizer10_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed11 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_304 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_305;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed12 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed12 <= main_mon_bussynchronizer11_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed12 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_305 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_306;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed13 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed13 <= main_mon_bussynchronizer12_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed13 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_306 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_307;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed14 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed14 <= main_mon_bussynchronizer13_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed14 <= main_mon_bussynchronizer14_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed14 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_307 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_308;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed15 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed15 <= main_mon_bussynchronizer15_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed15 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_308 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_309;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed16 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed16 <= main_mon_bussynchronizer16_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed16 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_309 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_310;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed17 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed17 <= main_mon_bussynchronizer17_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed17 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_310 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_311;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed18 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed18 <= main_mon_bussynchronizer18_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed18 <= main_mon_bussynchronizer19_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed18 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_311 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_312;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed19 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed19 <= main_mon_bussynchronizer20_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed19 <= main_mon_bussynchronizer21_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed19 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_312 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_313;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed20 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed20 <= main_mon_bussynchronizer22_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed20 <= main_mon_bussynchronizer23_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed20 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_313 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_314;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed21 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed21 <= main_mon_bussynchronizer24_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed21 <= main_mon_bussynchronizer25_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed21 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_314 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_315;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed22 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed22 <= main_mon_bussynchronizer26_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed22 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_315 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_316;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed23 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed23 <= main_mon_bussynchronizer27_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed23 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_316 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_317;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed24 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed24 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_317 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_318;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed25 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed25 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_318 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_319;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed26 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed26 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_319 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_320;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed27 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed27 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_320 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_321;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed28 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed28 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_321 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_322;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed29 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed29 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_322 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_323;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed30 <= 32'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer28_o;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer29_o;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer30_o;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer31_o;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer32_o;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer33_o;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer34_o;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer35_o;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer36_o;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer37_o;
		end
		default: begin
			builder_sync_t_rhs_array_muxed30 <= main_mon_bussynchronizer38_o;
		end
	endcase
// synthesis translate_off
	dummy_d_323 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_324;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed31 <= 1'd0;
	case (main_mon_probe_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
		default: begin
			builder_sync_t_rhs_array_muxed31 <= 1'd0;
		end
	endcase
// synthesis translate_off
	dummy_d_324 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_325;
// synthesis translate_on
always @(*) begin
	builder_sync_t_rhs_array_muxed2 <= 32'd0;
	case (main_mon_chan_sel_storage)
		1'd0: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed3;
		end
		1'd1: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed4;
		end
		2'd2: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed5;
		end
		2'd3: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed6;
		end
		3'd4: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed7;
		end
		3'd5: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed8;
		end
		3'd6: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed9;
		end
		3'd7: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed10;
		end
		4'd8: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed11;
		end
		4'd9: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed12;
		end
		4'd10: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed13;
		end
		4'd11: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed14;
		end
		4'd12: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed15;
		end
		4'd13: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed16;
		end
		4'd14: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed17;
		end
		4'd15: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed18;
		end
		5'd16: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed19;
		end
		5'd17: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed20;
		end
		5'd18: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed21;
		end
		5'd19: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed22;
		end
		5'd20: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed23;
		end
		5'd21: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed24;
		end
		5'd22: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed25;
		end
		5'd23: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed26;
		end
		5'd24: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed27;
		end
		5'd25: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed28;
		end
		5'd26: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed29;
		end
		5'd27: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed30;
		end
		default: begin
			builder_sync_t_rhs_array_muxed2 <= builder_sync_t_rhs_array_muxed31;
		end
	endcase
// synthesis translate_off
	dummy_d_325 <= dummy_s;
// synthesis translate_on
end
assign main_nist_clock_nist_clock_uart_phy_rx = builder_xilinxmultiregimpl0_regs1;
assign builder_xilinxasyncresetsynchronizerimpl0 = ((~main_nist_clock_pll_locked) | cpu_reset);
assign builder_xilinxasyncresetsynchronizerimpl1 = ((~main_nist_clock_pll_locked) | cpu_reset);
assign main_ethphy_toggle_o = builder_xilinxmultiregimpl1_regs1;
assign main_ps_preamble_error_toggle_o = builder_xilinxmultiregimpl2_regs1;
assign main_ps_crc_error_toggle_o = builder_xilinxmultiregimpl3_regs1;
assign main_tx_cdc_produce_rdomain = builder_xilinxmultiregimpl4_regs1;
assign main_tx_cdc_consume_wdomain = builder_xilinxmultiregimpl5_regs1;
assign main_rx_cdc_produce_rdomain = builder_xilinxmultiregimpl6_regs1;
assign main_rx_cdc_consume_wdomain = builder_xilinxmultiregimpl7_regs1;
assign main_i2c_status1 = builder_xilinxmultiregimpl8_regs1;
assign main_i2c_status2 = builder_xilinxmultiregimpl9_regs1;
assign builder_xilinxasyncresetsynchronizerimpl4 = (~main_rtio_crg_pll_locked);
assign main_rtio_crg_pll_locked_status = builder_xilinxmultiregimpl10_regs1;
assign main_value_gray_sys = builder_xilinxmultiregimpl11_regs1;
assign main_rtio_core_outputs_asyncfifobuffered0_produce_rdomain = builder_xilinxmultiregimpl12_regs1;
assign main_rtio_core_outputs_asyncfifobuffered0_consume_wdomain = builder_xilinxmultiregimpl13_regs1;
assign main_rtio_core_outputs_asyncfifobuffered1_produce_rdomain = builder_xilinxmultiregimpl14_regs1;
assign main_rtio_core_outputs_asyncfifobuffered1_consume_wdomain = builder_xilinxmultiregimpl15_regs1;
assign main_rtio_core_outputs_asyncfifobuffered2_produce_rdomain = builder_xilinxmultiregimpl16_regs1;
assign main_rtio_core_outputs_asyncfifobuffered2_consume_wdomain = builder_xilinxmultiregimpl17_regs1;
assign main_rtio_core_outputs_asyncfifobuffered3_produce_rdomain = builder_xilinxmultiregimpl18_regs1;
assign main_rtio_core_outputs_asyncfifobuffered3_consume_wdomain = builder_xilinxmultiregimpl19_regs1;
assign main_rtio_core_outputs_asyncfifobuffered4_produce_rdomain = builder_xilinxmultiregimpl20_regs1;
assign main_rtio_core_outputs_asyncfifobuffered4_consume_wdomain = builder_xilinxmultiregimpl21_regs1;
assign main_rtio_core_outputs_asyncfifobuffered5_produce_rdomain = builder_xilinxmultiregimpl22_regs1;
assign main_rtio_core_outputs_asyncfifobuffered5_consume_wdomain = builder_xilinxmultiregimpl23_regs1;
assign main_rtio_core_outputs_asyncfifobuffered6_produce_rdomain = builder_xilinxmultiregimpl24_regs1;
assign main_rtio_core_outputs_asyncfifobuffered6_consume_wdomain = builder_xilinxmultiregimpl25_regs1;
assign main_rtio_core_outputs_asyncfifobuffered7_produce_rdomain = builder_xilinxmultiregimpl26_regs1;
assign main_rtio_core_outputs_asyncfifobuffered7_consume_wdomain = builder_xilinxmultiregimpl27_regs1;
assign main_rtio_core_inputs_asyncfifo0_produce_rdomain = builder_xilinxmultiregimpl28_regs1;
assign main_rtio_core_inputs_asyncfifo0_consume_wdomain = builder_xilinxmultiregimpl29_regs1;
assign main_rtio_core_inputs_blindtransfer0_ps_toggle_o = builder_xilinxmultiregimpl30_regs1;
assign main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o = builder_xilinxmultiregimpl31_regs1;
assign main_rtio_core_inputs_asyncfifo1_produce_rdomain = builder_xilinxmultiregimpl32_regs1;
assign main_rtio_core_inputs_asyncfifo1_consume_wdomain = builder_xilinxmultiregimpl33_regs1;
assign main_rtio_core_inputs_blindtransfer1_ps_toggle_o = builder_xilinxmultiregimpl34_regs1;
assign main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o = builder_xilinxmultiregimpl35_regs1;
assign main_rtio_core_inputs_asyncfifo2_produce_rdomain = builder_xilinxmultiregimpl36_regs1;
assign main_rtio_core_inputs_asyncfifo2_consume_wdomain = builder_xilinxmultiregimpl37_regs1;
assign main_rtio_core_inputs_blindtransfer2_ps_toggle_o = builder_xilinxmultiregimpl38_regs1;
assign main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o = builder_xilinxmultiregimpl39_regs1;
assign main_rtio_core_inputs_asyncfifo3_produce_rdomain = builder_xilinxmultiregimpl40_regs1;
assign main_rtio_core_inputs_asyncfifo3_consume_wdomain = builder_xilinxmultiregimpl41_regs1;
assign main_rtio_core_inputs_blindtransfer3_ps_toggle_o = builder_xilinxmultiregimpl42_regs1;
assign main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o = builder_xilinxmultiregimpl43_regs1;
assign main_rtio_core_inputs_asyncfifo4_produce_rdomain = builder_xilinxmultiregimpl44_regs1;
assign main_rtio_core_inputs_asyncfifo4_consume_wdomain = builder_xilinxmultiregimpl45_regs1;
assign main_rtio_core_inputs_blindtransfer4_ps_toggle_o = builder_xilinxmultiregimpl46_regs1;
assign main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o = builder_xilinxmultiregimpl47_regs1;
assign main_rtio_core_inputs_asyncfifo5_produce_rdomain = builder_xilinxmultiregimpl48_regs1;
assign main_rtio_core_inputs_asyncfifo5_consume_wdomain = builder_xilinxmultiregimpl49_regs1;
assign main_rtio_core_inputs_blindtransfer5_ps_toggle_o = builder_xilinxmultiregimpl50_regs1;
assign main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o = builder_xilinxmultiregimpl51_regs1;
assign main_rtio_core_inputs_asyncfifo6_produce_rdomain = builder_xilinxmultiregimpl52_regs1;
assign main_rtio_core_inputs_asyncfifo6_consume_wdomain = builder_xilinxmultiregimpl53_regs1;
assign main_rtio_core_inputs_blindtransfer6_ps_toggle_o = builder_xilinxmultiregimpl54_regs1;
assign main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o = builder_xilinxmultiregimpl55_regs1;
assign main_rtio_core_inputs_asyncfifo7_produce_rdomain = builder_xilinxmultiregimpl56_regs1;
assign main_rtio_core_inputs_asyncfifo7_consume_wdomain = builder_xilinxmultiregimpl57_regs1;
assign main_rtio_core_inputs_blindtransfer7_ps_toggle_o = builder_xilinxmultiregimpl58_regs1;
assign main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o = builder_xilinxmultiregimpl59_regs1;
assign main_rtio_core_inputs_asyncfifo8_produce_rdomain = builder_xilinxmultiregimpl60_regs1;
assign main_rtio_core_inputs_asyncfifo8_consume_wdomain = builder_xilinxmultiregimpl61_regs1;
assign main_rtio_core_inputs_blindtransfer8_ps_toggle_o = builder_xilinxmultiregimpl62_regs1;
assign main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o = builder_xilinxmultiregimpl63_regs1;
assign main_rtio_core_inputs_asyncfifo9_produce_rdomain = builder_xilinxmultiregimpl64_regs1;
assign main_rtio_core_inputs_asyncfifo9_consume_wdomain = builder_xilinxmultiregimpl65_regs1;
assign main_rtio_core_inputs_blindtransfer9_ps_toggle_o = builder_xilinxmultiregimpl66_regs1;
assign main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o = builder_xilinxmultiregimpl67_regs1;
assign main_rtio_core_inputs_asyncfifo10_produce_rdomain = builder_xilinxmultiregimpl68_regs1;
assign main_rtio_core_inputs_asyncfifo10_consume_wdomain = builder_xilinxmultiregimpl69_regs1;
assign main_rtio_core_inputs_blindtransfer10_ps_toggle_o = builder_xilinxmultiregimpl70_regs1;
assign main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o = builder_xilinxmultiregimpl71_regs1;
assign main_rtio_core_inputs_asyncfifo11_produce_rdomain = builder_xilinxmultiregimpl72_regs1;
assign main_rtio_core_inputs_asyncfifo11_consume_wdomain = builder_xilinxmultiregimpl73_regs1;
assign main_rtio_core_inputs_blindtransfer11_ps_toggle_o = builder_xilinxmultiregimpl74_regs1;
assign main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o = builder_xilinxmultiregimpl75_regs1;
assign main_rtio_core_o_collision_sync_ps_toggle_o = builder_xilinxmultiregimpl76_regs1;
assign main_rtio_core_o_collision_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl77_regs1;
assign main_rtio_core_o_collision_sync_data_o = builder_xilinxmultiregimpl78_regs1;
assign main_rtio_core_o_busy_sync_ps_toggle_o = builder_xilinxmultiregimpl79_regs1;
assign main_rtio_core_o_busy_sync_ps_ack_toggle_o = builder_xilinxmultiregimpl80_regs1;
assign main_rtio_core_o_busy_sync_data_o = builder_xilinxmultiregimpl81_regs1;
assign main_mon_bussynchronizer0_o = builder_xilinxmultiregimpl82_regs1;
assign main_mon_bussynchronizer1_o = builder_xilinxmultiregimpl83_regs1;
assign main_mon_bussynchronizer2_o = builder_xilinxmultiregimpl84_regs1;
assign main_mon_bussynchronizer3_o = builder_xilinxmultiregimpl85_regs1;
assign main_mon_bussynchronizer4_o = builder_xilinxmultiregimpl86_regs1;
assign main_mon_bussynchronizer5_o = builder_xilinxmultiregimpl87_regs1;
assign main_mon_bussynchronizer6_o = builder_xilinxmultiregimpl88_regs1;
assign main_mon_bussynchronizer7_o = builder_xilinxmultiregimpl89_regs1;
assign main_mon_bussynchronizer8_o = builder_xilinxmultiregimpl90_regs1;
assign main_mon_bussynchronizer9_o = builder_xilinxmultiregimpl91_regs1;
assign main_mon_bussynchronizer10_o = builder_xilinxmultiregimpl92_regs1;
assign main_mon_bussynchronizer11_o = builder_xilinxmultiregimpl93_regs1;
assign main_mon_bussynchronizer12_o = builder_xilinxmultiregimpl94_regs1;
assign main_mon_bussynchronizer13_o = builder_xilinxmultiregimpl95_regs1;
assign main_mon_bussynchronizer14_o = builder_xilinxmultiregimpl96_regs1;
assign main_mon_bussynchronizer15_o = builder_xilinxmultiregimpl97_regs1;
assign main_mon_bussynchronizer16_o = builder_xilinxmultiregimpl98_regs1;
assign main_mon_bussynchronizer17_o = builder_xilinxmultiregimpl99_regs1;
assign main_mon_bussynchronizer18_o = builder_xilinxmultiregimpl100_regs1;
assign main_mon_bussynchronizer19_o = builder_xilinxmultiregimpl101_regs1;
assign main_mon_bussynchronizer20_o = builder_xilinxmultiregimpl102_regs1;
assign main_mon_bussynchronizer21_o = builder_xilinxmultiregimpl103_regs1;
assign main_mon_bussynchronizer22_o = builder_xilinxmultiregimpl104_regs1;
assign main_mon_bussynchronizer23_o = builder_xilinxmultiregimpl105_regs1;
assign main_mon_bussynchronizer24_o = builder_xilinxmultiregimpl106_regs1;
assign main_mon_bussynchronizer25_o = builder_xilinxmultiregimpl107_regs1;
assign main_mon_bussynchronizer26_o = builder_xilinxmultiregimpl108_regs1;
assign main_mon_bussynchronizer27_o = builder_xilinxmultiregimpl109_regs1;
assign main_mon_bussynchronizer28_ping_toggle_o = builder_xilinxmultiregimpl110_regs1;
assign main_mon_bussynchronizer28_pong_toggle_o = builder_xilinxmultiregimpl111_regs1;
assign main_mon_bussynchronizer28_obuffer = builder_xilinxmultiregimpl112_regs1;
assign main_mon_bussynchronizer29_ping_toggle_o = builder_xilinxmultiregimpl113_regs1;
assign main_mon_bussynchronizer29_pong_toggle_o = builder_xilinxmultiregimpl114_regs1;
assign main_mon_bussynchronizer29_obuffer = builder_xilinxmultiregimpl115_regs1;
assign main_mon_bussynchronizer30_ping_toggle_o = builder_xilinxmultiregimpl116_regs1;
assign main_mon_bussynchronizer30_pong_toggle_o = builder_xilinxmultiregimpl117_regs1;
assign main_mon_bussynchronizer30_obuffer = builder_xilinxmultiregimpl118_regs1;
assign main_mon_bussynchronizer31_ping_toggle_o = builder_xilinxmultiregimpl119_regs1;
assign main_mon_bussynchronizer31_pong_toggle_o = builder_xilinxmultiregimpl120_regs1;
assign main_mon_bussynchronizer31_obuffer = builder_xilinxmultiregimpl121_regs1;
assign main_mon_bussynchronizer32_ping_toggle_o = builder_xilinxmultiregimpl122_regs1;
assign main_mon_bussynchronizer32_pong_toggle_o = builder_xilinxmultiregimpl123_regs1;
assign main_mon_bussynchronizer32_obuffer = builder_xilinxmultiregimpl124_regs1;
assign main_mon_bussynchronizer33_ping_toggle_o = builder_xilinxmultiregimpl125_regs1;
assign main_mon_bussynchronizer33_pong_toggle_o = builder_xilinxmultiregimpl126_regs1;
assign main_mon_bussynchronizer33_obuffer = builder_xilinxmultiregimpl127_regs1;
assign main_mon_bussynchronizer34_ping_toggle_o = builder_xilinxmultiregimpl128_regs1;
assign main_mon_bussynchronizer34_pong_toggle_o = builder_xilinxmultiregimpl129_regs1;
assign main_mon_bussynchronizer34_obuffer = builder_xilinxmultiregimpl130_regs1;
assign main_mon_bussynchronizer35_ping_toggle_o = builder_xilinxmultiregimpl131_regs1;
assign main_mon_bussynchronizer35_pong_toggle_o = builder_xilinxmultiregimpl132_regs1;
assign main_mon_bussynchronizer35_obuffer = builder_xilinxmultiregimpl133_regs1;
assign main_mon_bussynchronizer36_ping_toggle_o = builder_xilinxmultiregimpl134_regs1;
assign main_mon_bussynchronizer36_pong_toggle_o = builder_xilinxmultiregimpl135_regs1;
assign main_mon_bussynchronizer36_obuffer = builder_xilinxmultiregimpl136_regs1;
assign main_mon_bussynchronizer37_ping_toggle_o = builder_xilinxmultiregimpl137_regs1;
assign main_mon_bussynchronizer37_pong_toggle_o = builder_xilinxmultiregimpl138_regs1;
assign main_mon_bussynchronizer37_obuffer = builder_xilinxmultiregimpl139_regs1;
assign main_mon_bussynchronizer38_ping_toggle_o = builder_xilinxmultiregimpl140_regs1;
assign main_mon_bussynchronizer38_pong_toggle_o = builder_xilinxmultiregimpl141_regs1;
assign main_mon_bussynchronizer38_obuffer = builder_xilinxmultiregimpl142_regs1;
assign main_output_8x0_override_en = builder_xilinxmultiregimpl143_regs1;
assign main_output_8x0_override_o = builder_xilinxmultiregimpl144_regs1;
assign main_output_8x1_override_en = builder_xilinxmultiregimpl145_regs1;
assign main_output_8x1_override_o = builder_xilinxmultiregimpl146_regs1;
assign main_output_8x2_override_en = builder_xilinxmultiregimpl147_regs1;
assign main_output_8x2_override_o = builder_xilinxmultiregimpl148_regs1;
assign main_inout_8x0_inout_8x0_override_en = builder_xilinxmultiregimpl149_regs1;
assign main_inout_8x0_inout_8x0_override_o = builder_xilinxmultiregimpl150_regs1;
assign main_inout_8x0_inout_8x0_override_oe = builder_xilinxmultiregimpl151_regs1;
assign main_output_8x3_override_en = builder_xilinxmultiregimpl152_regs1;
assign main_output_8x3_override_o = builder_xilinxmultiregimpl153_regs1;
assign main_output_8x4_override_en = builder_xilinxmultiregimpl154_regs1;
assign main_output_8x4_override_o = builder_xilinxmultiregimpl155_regs1;
assign main_output_8x5_override_en = builder_xilinxmultiregimpl156_regs1;
assign main_output_8x5_override_o = builder_xilinxmultiregimpl157_regs1;
assign main_inout_8x1_inout_8x1_override_en = builder_xilinxmultiregimpl158_regs1;
assign main_inout_8x1_inout_8x1_override_o = builder_xilinxmultiregimpl159_regs1;
assign main_inout_8x1_inout_8x1_override_oe = builder_xilinxmultiregimpl160_regs1;
assign main_output_8x6_override_en = builder_xilinxmultiregimpl161_regs1;
assign main_output_8x6_override_o = builder_xilinxmultiregimpl162_regs1;
assign main_output_8x7_override_en = builder_xilinxmultiregimpl163_regs1;
assign main_output_8x7_override_o = builder_xilinxmultiregimpl164_regs1;
assign main_output_8x8_override_en = builder_xilinxmultiregimpl165_regs1;
assign main_output_8x8_override_o = builder_xilinxmultiregimpl166_regs1;
assign main_inout_8x2_inout_8x2_override_en = builder_xilinxmultiregimpl167_regs1;
assign main_inout_8x2_inout_8x2_override_o = builder_xilinxmultiregimpl168_regs1;
assign main_inout_8x2_inout_8x2_override_oe = builder_xilinxmultiregimpl169_regs1;
assign main_output_8x9_override_en = builder_xilinxmultiregimpl170_regs1;
assign main_output_8x9_override_o = builder_xilinxmultiregimpl171_regs1;
assign main_output_8x10_override_en = builder_xilinxmultiregimpl172_regs1;
assign main_output_8x10_override_o = builder_xilinxmultiregimpl173_regs1;
assign main_output_8x11_override_en = builder_xilinxmultiregimpl174_regs1;
assign main_output_8x11_override_o = builder_xilinxmultiregimpl175_regs1;
assign main_inout_8x3_inout_8x3_override_en = builder_xilinxmultiregimpl176_regs1;
assign main_inout_8x3_inout_8x3_override_o = builder_xilinxmultiregimpl177_regs1;
assign main_inout_8x3_inout_8x3_override_oe = builder_xilinxmultiregimpl178_regs1;
assign main_inout_8x4_inout_8x4_override_en = builder_xilinxmultiregimpl179_regs1;
assign main_inout_8x4_inout_8x4_override_o = builder_xilinxmultiregimpl180_regs1;
assign main_inout_8x4_inout_8x4_override_oe = builder_xilinxmultiregimpl181_regs1;
assign main_inout_8x5_inout_8x5_override_en = builder_xilinxmultiregimpl182_regs1;
assign main_inout_8x5_inout_8x5_override_o = builder_xilinxmultiregimpl183_regs1;
assign main_inout_8x5_inout_8x5_override_oe = builder_xilinxmultiregimpl184_regs1;
assign main_inout_8x6_inout_8x6_override_en = builder_xilinxmultiregimpl185_regs1;
assign main_inout_8x6_inout_8x6_override_o = builder_xilinxmultiregimpl186_regs1;
assign main_inout_8x6_inout_8x6_override_oe = builder_xilinxmultiregimpl187_regs1;
assign main_output0_override_en = builder_xilinxmultiregimpl188_regs1;
assign main_output0_override_o = builder_xilinxmultiregimpl189_regs1;
assign main_output1_override_en = builder_xilinxmultiregimpl190_regs1;
assign main_output1_override_o = builder_xilinxmultiregimpl191_regs1;

always @(posedge clk200_clk) begin
	if ((main_nist_clock_reset_counter != 1'd0)) begin
		main_nist_clock_reset_counter <= (main_nist_clock_reset_counter - 1'd1);
	end else begin
		main_nist_clock_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		main_nist_clock_reset_counter <= 4'd15;
		main_nist_clock_ic_reset <= 1'd1;
	end
end

always @(posedge eth_rx_clk) begin
	main_ethphy_eth_counter <= (main_ethphy_eth_counter + 1'd1);
	if (main_ethphy_i) begin
		main_ethphy_toggle_i <= (~main_ethphy_toggle_i);
	end
	main_ethphy_liteethphygmiimiirx_pads_d_rx_dv <= eth_rx_dv;
	main_ethphy_liteethphygmiimiirx_pads_d_rx_data <= eth_rx_data;
	main_ethphy_liteethphygmiimiirx_gmii_rx_rx_dv_d <= main_ethphy_liteethphygmiimiirx_pads_d_rx_dv;
	main_ethphy_liteethphygmiimiirx_gmii_rx_source_stb <= main_ethphy_liteethphygmiimiirx_pads_d_rx_dv;
	main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_data <= main_ethphy_liteethphygmiimiirx_pads_d_rx_data;
	main_ethphy_liteethphygmiimiirx_converter_reset <= (~main_ethphy_liteethphygmiimiirx_pads_d_rx_dv);
	main_ethphy_liteethphygmiimiirx_converter_sink_stb <= 1'd1;
	main_ethphy_liteethphygmiimiirx_converter_sink_payload_data <= main_ethphy_liteethphygmiimiirx_pads_d_rx_data;
	if (main_ethphy_liteethphygmiimiirx_converter_source_ack) begin
		main_ethphy_liteethphygmiimiirx_converter_strobe_all <= 1'd0;
	end
	if (main_ethphy_liteethphygmiimiirx_converter_load_part) begin
		if (((main_ethphy_liteethphygmiimiirx_converter_demux == 1'd1) | main_ethphy_liteethphygmiimiirx_converter_sink_eop)) begin
			main_ethphy_liteethphygmiimiirx_converter_demux <= 1'd0;
			main_ethphy_liteethphygmiimiirx_converter_strobe_all <= 1'd1;
		end else begin
			main_ethphy_liteethphygmiimiirx_converter_demux <= (main_ethphy_liteethphygmiimiirx_converter_demux + 1'd1);
		end
	end
	if ((main_ethphy_liteethphygmiimiirx_converter_source_stb & main_ethphy_liteethphygmiimiirx_converter_source_ack)) begin
		main_ethphy_liteethphygmiimiirx_converter_source_eop <= main_ethphy_liteethphygmiimiirx_converter_sink_eop;
	end else begin
		if ((main_ethphy_liteethphygmiimiirx_converter_sink_stb & main_ethphy_liteethphygmiimiirx_converter_sink_ack)) begin
			main_ethphy_liteethphygmiimiirx_converter_source_eop <= (main_ethphy_liteethphygmiimiirx_converter_sink_eop | main_ethphy_liteethphygmiimiirx_converter_source_eop);
		end
	end
	if (main_ethphy_liteethphygmiimiirx_converter_load_part) begin
		case (main_ethphy_liteethphygmiimiirx_converter_demux)
			1'd0: begin
				main_ethphy_liteethphygmiimiirx_converter_source_payload_data[3:0] <= main_ethphy_liteethphygmiimiirx_converter_sink_payload_data;
			end
			1'd1: begin
				main_ethphy_liteethphygmiimiirx_converter_source_payload_data[7:4] <= main_ethphy_liteethphygmiimiirx_converter_sink_payload_data;
			end
		endcase
	end
	if (main_ethphy_liteethphygmiimiirx_converter_reset) begin
		main_ethphy_liteethphygmiimiirx_converter_source_eop <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_source_payload_data <= 8'd0;
		main_ethphy_liteethphygmiimiirx_converter_demux <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_strobe_all <= 1'd0;
	end
	builder_liteethmacpreamblechecker_state <= builder_liteethmacpreamblechecker_next_state;
	if (main_crc32_checker_crc_ce) begin
		main_crc32_checker_crc_reg <= main_crc32_checker_crc_next;
	end
	if (main_crc32_checker_crc_reset) begin
		main_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((main_crc32_checker_syncfifo_syncfifo_we & main_crc32_checker_syncfifo_syncfifo_writable) & (~main_crc32_checker_syncfifo_replace))) begin
		if ((main_crc32_checker_syncfifo_produce == 3'd4)) begin
			main_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			main_crc32_checker_syncfifo_produce <= (main_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (main_crc32_checker_syncfifo_do_read) begin
		if ((main_crc32_checker_syncfifo_consume == 3'd4)) begin
			main_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			main_crc32_checker_syncfifo_consume <= (main_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((main_crc32_checker_syncfifo_syncfifo_we & main_crc32_checker_syncfifo_syncfifo_writable) & (~main_crc32_checker_syncfifo_replace))) begin
		if ((~main_crc32_checker_syncfifo_do_read)) begin
			main_crc32_checker_syncfifo_level <= (main_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (main_crc32_checker_syncfifo_do_read) begin
			main_crc32_checker_syncfifo_level <= (main_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (main_crc32_checker_fifo_reset) begin
		main_crc32_checker_syncfifo_level <= 3'd0;
		main_crc32_checker_syncfifo_produce <= 3'd0;
		main_crc32_checker_syncfifo_consume <= 3'd0;
	end
	builder_liteethmaccrc32checker_state <= builder_liteethmaccrc32checker_next_state;
	if (main_ps_preamble_error_i) begin
		main_ps_preamble_error_toggle_i <= (~main_ps_preamble_error_toggle_i);
	end
	if (main_ps_crc_error_i) begin
		main_ps_crc_error_toggle_i <= (~main_ps_crc_error_toggle_i);
	end
	if (main_rx_converter_converter_source_ack) begin
		main_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (main_rx_converter_converter_load_part) begin
		if (((main_rx_converter_converter_demux == 2'd3) | main_rx_converter_converter_sink_eop)) begin
			main_rx_converter_converter_demux <= 1'd0;
			main_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			main_rx_converter_converter_demux <= (main_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((main_rx_converter_converter_source_stb & main_rx_converter_converter_source_ack)) begin
		main_rx_converter_converter_source_eop <= main_rx_converter_converter_sink_eop;
	end else begin
		if ((main_rx_converter_converter_sink_stb & main_rx_converter_converter_sink_ack)) begin
			main_rx_converter_converter_source_eop <= (main_rx_converter_converter_sink_eop | main_rx_converter_converter_source_eop);
		end
	end
	if (main_rx_converter_converter_load_part) begin
		case (main_rx_converter_converter_demux)
			1'd0: begin
				main_rx_converter_converter_source_payload_data[39:30] <= main_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				main_rx_converter_converter_source_payload_data[29:20] <= main_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				main_rx_converter_converter_source_payload_data[19:10] <= main_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				main_rx_converter_converter_source_payload_data[9:0] <= main_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	main_rx_cdc_graycounter0_q_binary <= main_rx_cdc_graycounter0_q_next_binary;
	main_rx_cdc_graycounter0_q <= main_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		main_ethphy_eth_counter <= 10'd0;
		main_ethphy_liteethphygmiimiirx_pads_d_rx_dv <= 1'd0;
		main_ethphy_liteethphygmiimiirx_pads_d_rx_data <= 8'd0;
		main_ethphy_liteethphygmiimiirx_gmii_rx_source_stb <= 1'd0;
		main_ethphy_liteethphygmiimiirx_gmii_rx_source_payload_data <= 8'd0;
		main_ethphy_liteethphygmiimiirx_gmii_rx_rx_dv_d <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_sink_stb <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_sink_payload_data <= 4'd0;
		main_ethphy_liteethphygmiimiirx_converter_source_eop <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_source_payload_data <= 8'd0;
		main_ethphy_liteethphygmiimiirx_converter_demux <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_strobe_all <= 1'd0;
		main_ethphy_liteethphygmiimiirx_converter_reset <= 1'd0;
		main_crc32_checker_crc_reg <= 32'd4294967295;
		main_crc32_checker_syncfifo_level <= 3'd0;
		main_crc32_checker_syncfifo_produce <= 3'd0;
		main_crc32_checker_syncfifo_consume <= 3'd0;
		main_rx_converter_converter_source_eop <= 1'd0;
		main_rx_converter_converter_source_payload_data <= 40'd0;
		main_rx_converter_converter_demux <= 2'd0;
		main_rx_converter_converter_strobe_all <= 1'd0;
		main_rx_cdc_graycounter0_q <= 7'd0;
		main_rx_cdc_graycounter0_q_binary <= 7'd0;
		builder_liteethmacpreamblechecker_state <= 1'd0;
		builder_liteethmaccrc32checker_state <= 2'd0;
	end
	builder_xilinxmultiregimpl7_regs0 <= main_rx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl7_regs1 <= builder_xilinxmultiregimpl7_regs0;
end

always @(posedge eth_tx_clk) begin
	if ((main_ethphy_mode0 == 1'd1)) begin
		eth_tx_en <= main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_en;
		eth_tx_data <= main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_data;
	end else begin
		eth_tx_en <= main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_en;
		eth_tx_data <= main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_data;
	end
	main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_er <= 1'd0;
	main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_en <= main_ethphy_liteethphygmiimiitx_gmii_tx_sink_stb;
	main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_data <= main_ethphy_liteethphygmiimiitx_gmii_tx_sink_payload_data;
	main_ethphy_liteethphygmiimiitx_gmii_tx_sink_ack <= 1'd1;
	main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_er <= 1'd0;
	main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_en <= main_ethphy_liteethphygmiimiitx_converter_source_stb;
	main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_data <= main_ethphy_liteethphygmiimiitx_converter_source_payload_data;
	if ((main_ethphy_liteethphygmiimiitx_converter_source_stb & main_ethphy_liteethphygmiimiitx_converter_source_ack)) begin
		if (main_ethphy_liteethphygmiimiitx_converter_last) begin
			main_ethphy_liteethphygmiimiitx_converter_mux <= 1'd0;
		end else begin
			main_ethphy_liteethphygmiimiitx_converter_mux <= (main_ethphy_liteethphygmiimiitx_converter_mux + 1'd1);
		end
	end
	if (main_tx_gap_inserter_counter_reset) begin
		main_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (main_tx_gap_inserter_counter_ce) begin
			main_tx_gap_inserter_counter <= (main_tx_gap_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacgap_state <= builder_liteethmacgap_next_state;
	if (main_preamble_inserter_clr_cnt) begin
		main_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (main_preamble_inserter_inc_cnt) begin
			main_preamble_inserter_cnt <= (main_preamble_inserter_cnt + 1'd1);
		end
	end
	builder_liteethmacpreambleinserter_state <= builder_liteethmacpreambleinserter_next_state;
	if (main_crc32_inserter_is_ongoing0) begin
		main_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((main_crc32_inserter_is_ongoing1 & (~main_crc32_inserter_cnt_done))) begin
			main_crc32_inserter_cnt <= (main_crc32_inserter_cnt - main_crc32_inserter_source_ack);
		end
	end
	if (main_crc32_inserter_ce) begin
		main_crc32_inserter_reg <= main_crc32_inserter_next;
	end
	if (main_crc32_inserter_reset) begin
		main_crc32_inserter_reg <= 32'd4294967295;
	end
	builder_liteethmaccrc32inserter_state <= builder_liteethmaccrc32inserter_next_state;
	if (main_padding_inserter_counter_reset) begin
		main_padding_inserter_counter <= 1'd0;
	end else begin
		if (main_padding_inserter_counter_ce) begin
			main_padding_inserter_counter <= (main_padding_inserter_counter + 1'd1);
		end
	end
	builder_liteethmacpaddinginserter_state <= builder_liteethmacpaddinginserter_next_state;
	if ((main_tx_last_be_sink_stb & main_tx_last_be_sink_ack)) begin
		if (main_tx_last_be_sink_eop) begin
			main_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (main_tx_last_be_sink_payload_last_be) begin
				main_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((main_tx_converter_converter_source_stb & main_tx_converter_converter_source_ack)) begin
		if (main_tx_converter_converter_last) begin
			main_tx_converter_converter_mux <= 1'd0;
		end else begin
			main_tx_converter_converter_mux <= (main_tx_converter_converter_mux + 1'd1);
		end
	end
	main_tx_cdc_graycounter1_q_binary <= main_tx_cdc_graycounter1_q_next_binary;
	main_tx_cdc_graycounter1_q <= main_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		eth_tx_en <= 1'd0;
		eth_tx_data <= 8'd0;
		main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_er <= 1'd0;
		main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_en <= 1'd0;
		main_ethphy_liteethphygmiimiitx_gmii_tx_pads_tx_data <= 8'd0;
		main_ethphy_liteethphygmiimiitx_gmii_tx_sink_ack <= 1'd0;
		main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_er <= 1'd0;
		main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_en <= 1'd0;
		main_ethphy_liteethphygmiimiitx_mii_tx_pads_tx_data <= 8'd0;
		main_ethphy_liteethphygmiimiitx_converter_mux <= 1'd0;
		main_tx_gap_inserter_counter <= 4'd0;
		main_preamble_inserter_cnt <= 3'd0;
		main_crc32_inserter_reg <= 32'd4294967295;
		main_crc32_inserter_cnt <= 2'd3;
		main_padding_inserter_counter <= 16'd1;
		main_tx_last_be_ongoing <= 1'd1;
		main_tx_converter_converter_mux <= 2'd0;
		main_tx_cdc_graycounter1_q <= 7'd0;
		main_tx_cdc_graycounter1_q_binary <= 7'd0;
		builder_liteethmacgap_state <= 1'd0;
		builder_liteethmacpreambleinserter_state <= 2'd0;
		builder_liteethmaccrc32inserter_state <= 2'd0;
		builder_liteethmacpaddinginserter_state <= 1'd0;
	end
	builder_xilinxmultiregimpl4_regs0 <= main_tx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl4_regs1 <= builder_xilinxmultiregimpl4_regs0;
end

always @(posedge ext_clkout_clk) begin
	user_sma_gpio_p_33 <= (~user_sma_gpio_p_33);
end

always @(posedge rio_clk) begin
	main_inout_8x0_inout_8x0_sample <= 1'd0;
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & main_inout_8x0_inout_8x0_ointerface0_address[1])) begin
		main_inout_8x0_inout_8x0_sensitivity <= main_inout_8x0_inout_8x0_ointerface0_data;
		if (main_inout_8x0_inout_8x0_ointerface0_address[0]) begin
			main_inout_8x0_inout_8x0_sample <= 1'd1;
		end
	end
	main_inout_8x1_inout_8x1_sample <= 1'd0;
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & main_inout_8x1_inout_8x1_ointerface1_address[1])) begin
		main_inout_8x1_inout_8x1_sensitivity <= main_inout_8x1_inout_8x1_ointerface1_data;
		if (main_inout_8x1_inout_8x1_ointerface1_address[0]) begin
			main_inout_8x1_inout_8x1_sample <= 1'd1;
		end
	end
	main_inout_8x2_inout_8x2_sample <= 1'd0;
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & main_inout_8x2_inout_8x2_ointerface2_address[1])) begin
		main_inout_8x2_inout_8x2_sensitivity <= main_inout_8x2_inout_8x2_ointerface2_data;
		if (main_inout_8x2_inout_8x2_ointerface2_address[0]) begin
			main_inout_8x2_inout_8x2_sample <= 1'd1;
		end
	end
	main_inout_8x3_inout_8x3_sample <= 1'd0;
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & main_inout_8x3_inout_8x3_ointerface3_address[1])) begin
		main_inout_8x3_inout_8x3_sensitivity <= main_inout_8x3_inout_8x3_ointerface3_data;
		if (main_inout_8x3_inout_8x3_ointerface3_address[0]) begin
			main_inout_8x3_inout_8x3_sample <= 1'd1;
		end
	end
	main_inout_8x4_inout_8x4_sample <= 1'd0;
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & main_inout_8x4_inout_8x4_ointerface4_address[1])) begin
		main_inout_8x4_inout_8x4_sensitivity <= main_inout_8x4_inout_8x4_ointerface4_data;
		if (main_inout_8x4_inout_8x4_ointerface4_address[0]) begin
			main_inout_8x4_inout_8x4_sample <= 1'd1;
		end
	end
	main_inout_8x5_inout_8x5_sample <= 1'd0;
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & main_inout_8x5_inout_8x5_ointerface5_address[1])) begin
		main_inout_8x5_inout_8x5_sensitivity <= main_inout_8x5_inout_8x5_ointerface5_data;
		if (main_inout_8x5_inout_8x5_ointerface5_address[0]) begin
			main_inout_8x5_inout_8x5_sample <= 1'd1;
		end
	end
	main_inout_8x6_inout_8x6_sample <= 1'd0;
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & main_inout_8x6_inout_8x6_ointerface6_address[1])) begin
		main_inout_8x6_inout_8x6_sensitivity <= main_inout_8x6_inout_8x6_ointerface6_data;
		if (main_inout_8x6_inout_8x6_ointerface6_address[0]) begin
			main_inout_8x6_inout_8x6_sample <= 1'd1;
		end
	end
	if (main_clockgen_stb) begin
		main_clockgen_ftw <= main_clockgen_data;
	end
	if (main_ad9914_stb) begin
		main_ad9914_current_address <= main_ad9914_address;
		main_ad9914_current_data <= main_ad9914_data;
	end
	if ((main_ad9914_current_address == 8'd129)) begin
		main_ad9914_current_sel <= main_ad9914_current_data[15:1];
	end
	if (main_ad9914_stb) begin
		main_ad9914_active <= 1'd1;
		main_ad9914_bus_adr <= main_ad9914_address[7:0];
		main_ad9914_bus_we <= 1'd1;
		main_ad9914_bus_dat_w <= main_ad9914_data;
		main_ad9914_bus_sel <= 2'd3;
	end
	if (main_ad9914_bus_ack) begin
		main_ad9914_active <= 1'd0;
	end
	if ((main_rtio_core_outputs_asyncfifobuffered0_re | (~main_rtio_core_outputs_asyncfifobuffered0_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered0_dout <= main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_dout;
		main_rtio_core_outputs_asyncfifobuffered0_readable <= main_rtio_core_outputs_asyncfifobuffered0_asyncfifo0_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered1_re | (~main_rtio_core_outputs_asyncfifobuffered1_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered1_dout <= main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_dout;
		main_rtio_core_outputs_asyncfifobuffered1_readable <= main_rtio_core_outputs_asyncfifobuffered1_asyncfifo1_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered2_re | (~main_rtio_core_outputs_asyncfifobuffered2_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered2_dout <= main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_dout;
		main_rtio_core_outputs_asyncfifobuffered2_readable <= main_rtio_core_outputs_asyncfifobuffered2_asyncfifo2_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered3_re | (~main_rtio_core_outputs_asyncfifobuffered3_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered3_dout <= main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_dout;
		main_rtio_core_outputs_asyncfifobuffered3_readable <= main_rtio_core_outputs_asyncfifobuffered3_asyncfifo3_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered4_re | (~main_rtio_core_outputs_asyncfifobuffered4_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered4_dout <= main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_dout;
		main_rtio_core_outputs_asyncfifobuffered4_readable <= main_rtio_core_outputs_asyncfifobuffered4_asyncfifo4_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered5_re | (~main_rtio_core_outputs_asyncfifobuffered5_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered5_dout <= main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_dout;
		main_rtio_core_outputs_asyncfifobuffered5_readable <= main_rtio_core_outputs_asyncfifobuffered5_asyncfifo5_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered6_re | (~main_rtio_core_outputs_asyncfifobuffered6_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered6_dout <= main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_dout;
		main_rtio_core_outputs_asyncfifobuffered6_readable <= main_rtio_core_outputs_asyncfifobuffered6_asyncfifo6_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_next;
	if ((main_rtio_core_outputs_asyncfifobuffered7_re | (~main_rtio_core_outputs_asyncfifobuffered7_readable))) begin
		main_rtio_core_outputs_asyncfifobuffered7_dout <= main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_dout;
		main_rtio_core_outputs_asyncfifobuffered7_readable <= main_rtio_core_outputs_asyncfifobuffered7_asyncfifo7_readable;
	end
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_next;
	main_rtio_core_outputs_gates_record0_payload_channel1 <= main_rtio_core_outputs_gates_record0_payload_channel0;
	main_rtio_core_outputs_gates_record0_payload_fine_ts <= main_rtio_core_outputs_gates_record0_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record0_payload_address1 <= main_rtio_core_outputs_gates_record0_payload_address0;
	main_rtio_core_outputs_gates_record0_payload_data1 <= main_rtio_core_outputs_gates_record0_payload_data0;
	main_rtio_core_outputs_gates_record0_seqn1 <= main_rtio_core_outputs_gates_record0_seqn0;
	main_rtio_core_outputs_gates_record0_valid <= (main_rtio_core_outputs_gates_record0_re & main_rtio_core_outputs_gates_record0_readable);
	main_rtio_core_outputs_gates_record1_payload_channel1 <= main_rtio_core_outputs_gates_record1_payload_channel0;
	main_rtio_core_outputs_gates_record1_payload_fine_ts <= main_rtio_core_outputs_gates_record1_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record1_payload_address1 <= main_rtio_core_outputs_gates_record1_payload_address0;
	main_rtio_core_outputs_gates_record1_payload_data1 <= main_rtio_core_outputs_gates_record1_payload_data0;
	main_rtio_core_outputs_gates_record1_seqn1 <= main_rtio_core_outputs_gates_record1_seqn0;
	main_rtio_core_outputs_gates_record1_valid <= (main_rtio_core_outputs_gates_record1_re & main_rtio_core_outputs_gates_record1_readable);
	main_rtio_core_outputs_gates_record2_payload_channel1 <= main_rtio_core_outputs_gates_record2_payload_channel0;
	main_rtio_core_outputs_gates_record2_payload_fine_ts <= main_rtio_core_outputs_gates_record2_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record2_payload_address1 <= main_rtio_core_outputs_gates_record2_payload_address0;
	main_rtio_core_outputs_gates_record2_payload_data1 <= main_rtio_core_outputs_gates_record2_payload_data0;
	main_rtio_core_outputs_gates_record2_seqn1 <= main_rtio_core_outputs_gates_record2_seqn0;
	main_rtio_core_outputs_gates_record2_valid <= (main_rtio_core_outputs_gates_record2_re & main_rtio_core_outputs_gates_record2_readable);
	main_rtio_core_outputs_gates_record3_payload_channel1 <= main_rtio_core_outputs_gates_record3_payload_channel0;
	main_rtio_core_outputs_gates_record3_payload_fine_ts <= main_rtio_core_outputs_gates_record3_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record3_payload_address1 <= main_rtio_core_outputs_gates_record3_payload_address0;
	main_rtio_core_outputs_gates_record3_payload_data1 <= main_rtio_core_outputs_gates_record3_payload_data0;
	main_rtio_core_outputs_gates_record3_seqn1 <= main_rtio_core_outputs_gates_record3_seqn0;
	main_rtio_core_outputs_gates_record3_valid <= (main_rtio_core_outputs_gates_record3_re & main_rtio_core_outputs_gates_record3_readable);
	main_rtio_core_outputs_gates_record4_payload_channel1 <= main_rtio_core_outputs_gates_record4_payload_channel0;
	main_rtio_core_outputs_gates_record4_payload_fine_ts <= main_rtio_core_outputs_gates_record4_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record4_payload_address1 <= main_rtio_core_outputs_gates_record4_payload_address0;
	main_rtio_core_outputs_gates_record4_payload_data1 <= main_rtio_core_outputs_gates_record4_payload_data0;
	main_rtio_core_outputs_gates_record4_seqn1 <= main_rtio_core_outputs_gates_record4_seqn0;
	main_rtio_core_outputs_gates_record4_valid <= (main_rtio_core_outputs_gates_record4_re & main_rtio_core_outputs_gates_record4_readable);
	main_rtio_core_outputs_gates_record5_payload_channel1 <= main_rtio_core_outputs_gates_record5_payload_channel0;
	main_rtio_core_outputs_gates_record5_payload_fine_ts <= main_rtio_core_outputs_gates_record5_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record5_payload_address1 <= main_rtio_core_outputs_gates_record5_payload_address0;
	main_rtio_core_outputs_gates_record5_payload_data1 <= main_rtio_core_outputs_gates_record5_payload_data0;
	main_rtio_core_outputs_gates_record5_seqn1 <= main_rtio_core_outputs_gates_record5_seqn0;
	main_rtio_core_outputs_gates_record5_valid <= (main_rtio_core_outputs_gates_record5_re & main_rtio_core_outputs_gates_record5_readable);
	main_rtio_core_outputs_gates_record6_payload_channel1 <= main_rtio_core_outputs_gates_record6_payload_channel0;
	main_rtio_core_outputs_gates_record6_payload_fine_ts <= main_rtio_core_outputs_gates_record6_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record6_payload_address1 <= main_rtio_core_outputs_gates_record6_payload_address0;
	main_rtio_core_outputs_gates_record6_payload_data1 <= main_rtio_core_outputs_gates_record6_payload_data0;
	main_rtio_core_outputs_gates_record6_seqn1 <= main_rtio_core_outputs_gates_record6_seqn0;
	main_rtio_core_outputs_gates_record6_valid <= (main_rtio_core_outputs_gates_record6_re & main_rtio_core_outputs_gates_record6_readable);
	main_rtio_core_outputs_gates_record7_payload_channel1 <= main_rtio_core_outputs_gates_record7_payload_channel0;
	main_rtio_core_outputs_gates_record7_payload_fine_ts <= main_rtio_core_outputs_gates_record7_payload_timestamp[2:0];
	main_rtio_core_outputs_gates_record7_payload_address1 <= main_rtio_core_outputs_gates_record7_payload_address0;
	main_rtio_core_outputs_gates_record7_payload_data1 <= main_rtio_core_outputs_gates_record7_payload_data0;
	main_rtio_core_outputs_gates_record7_seqn1 <= main_rtio_core_outputs_gates_record7_seqn0;
	main_rtio_core_outputs_gates_record7_valid <= (main_rtio_core_outputs_gates_record7_re & main_rtio_core_outputs_gates_record7_readable);
	main_rtio_core_outputs_record0_valid1 <= main_rtio_core_outputs_record40_rec_valid;
	main_rtio_core_outputs_record0_payload_channel3 <= main_rtio_core_outputs_record40_rec_payload_channel;
	main_rtio_core_outputs_record0_payload_fine_ts1 <= main_rtio_core_outputs_record40_rec_payload_fine_ts;
	main_rtio_core_outputs_record0_payload_address3 <= main_rtio_core_outputs_record40_rec_payload_address;
	main_rtio_core_outputs_record0_payload_data3 <= main_rtio_core_outputs_record40_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r0 <= main_rtio_core_outputs_record40_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r0 <= main_rtio_core_outputs_record40_rec_nondata_replace_occured;
	main_rtio_core_outputs_record1_valid1 <= main_rtio_core_outputs_record41_rec_valid;
	main_rtio_core_outputs_record1_payload_channel3 <= main_rtio_core_outputs_record41_rec_payload_channel;
	main_rtio_core_outputs_record1_payload_fine_ts1 <= main_rtio_core_outputs_record41_rec_payload_fine_ts;
	main_rtio_core_outputs_record1_payload_address3 <= main_rtio_core_outputs_record41_rec_payload_address;
	main_rtio_core_outputs_record1_payload_data3 <= main_rtio_core_outputs_record41_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r1 <= main_rtio_core_outputs_record41_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r1 <= main_rtio_core_outputs_record41_rec_nondata_replace_occured;
	main_rtio_core_outputs_record2_valid1 <= main_rtio_core_outputs_record42_rec_valid;
	main_rtio_core_outputs_record2_payload_channel3 <= main_rtio_core_outputs_record42_rec_payload_channel;
	main_rtio_core_outputs_record2_payload_fine_ts1 <= main_rtio_core_outputs_record42_rec_payload_fine_ts;
	main_rtio_core_outputs_record2_payload_address3 <= main_rtio_core_outputs_record42_rec_payload_address;
	main_rtio_core_outputs_record2_payload_data3 <= main_rtio_core_outputs_record42_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r2 <= main_rtio_core_outputs_record42_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r2 <= main_rtio_core_outputs_record42_rec_nondata_replace_occured;
	main_rtio_core_outputs_record3_valid1 <= main_rtio_core_outputs_record43_rec_valid;
	main_rtio_core_outputs_record3_payload_channel3 <= main_rtio_core_outputs_record43_rec_payload_channel;
	main_rtio_core_outputs_record3_payload_fine_ts1 <= main_rtio_core_outputs_record43_rec_payload_fine_ts;
	main_rtio_core_outputs_record3_payload_address3 <= main_rtio_core_outputs_record43_rec_payload_address;
	main_rtio_core_outputs_record3_payload_data3 <= main_rtio_core_outputs_record43_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r3 <= main_rtio_core_outputs_record43_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r3 <= main_rtio_core_outputs_record43_rec_nondata_replace_occured;
	main_rtio_core_outputs_record4_valid1 <= main_rtio_core_outputs_record44_rec_valid;
	main_rtio_core_outputs_record4_payload_channel3 <= main_rtio_core_outputs_record44_rec_payload_channel;
	main_rtio_core_outputs_record4_payload_fine_ts1 <= main_rtio_core_outputs_record44_rec_payload_fine_ts;
	main_rtio_core_outputs_record4_payload_address3 <= main_rtio_core_outputs_record44_rec_payload_address;
	main_rtio_core_outputs_record4_payload_data3 <= main_rtio_core_outputs_record44_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r4 <= main_rtio_core_outputs_record44_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r4 <= main_rtio_core_outputs_record44_rec_nondata_replace_occured;
	main_rtio_core_outputs_record5_valid1 <= main_rtio_core_outputs_record45_rec_valid;
	main_rtio_core_outputs_record5_payload_channel3 <= main_rtio_core_outputs_record45_rec_payload_channel;
	main_rtio_core_outputs_record5_payload_fine_ts1 <= main_rtio_core_outputs_record45_rec_payload_fine_ts;
	main_rtio_core_outputs_record5_payload_address3 <= main_rtio_core_outputs_record45_rec_payload_address;
	main_rtio_core_outputs_record5_payload_data3 <= main_rtio_core_outputs_record45_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r5 <= main_rtio_core_outputs_record45_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r5 <= main_rtio_core_outputs_record45_rec_nondata_replace_occured;
	main_rtio_core_outputs_record6_valid1 <= main_rtio_core_outputs_record46_rec_valid;
	main_rtio_core_outputs_record6_payload_channel3 <= main_rtio_core_outputs_record46_rec_payload_channel;
	main_rtio_core_outputs_record6_payload_fine_ts1 <= main_rtio_core_outputs_record46_rec_payload_fine_ts;
	main_rtio_core_outputs_record6_payload_address3 <= main_rtio_core_outputs_record46_rec_payload_address;
	main_rtio_core_outputs_record6_payload_data3 <= main_rtio_core_outputs_record46_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r6 <= main_rtio_core_outputs_record46_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r6 <= main_rtio_core_outputs_record46_rec_nondata_replace_occured;
	main_rtio_core_outputs_record7_valid1 <= main_rtio_core_outputs_record47_rec_valid;
	main_rtio_core_outputs_record7_payload_channel3 <= main_rtio_core_outputs_record47_rec_payload_channel;
	main_rtio_core_outputs_record7_payload_fine_ts1 <= main_rtio_core_outputs_record47_rec_payload_fine_ts;
	main_rtio_core_outputs_record7_payload_address3 <= main_rtio_core_outputs_record47_rec_payload_address;
	main_rtio_core_outputs_record7_payload_data3 <= main_rtio_core_outputs_record47_rec_payload_data;
	main_rtio_core_outputs_replace_occured_r7 <= main_rtio_core_outputs_record47_rec_replace_occured;
	main_rtio_core_outputs_nondata_replace_occured_r7 <= main_rtio_core_outputs_record47_rec_nondata_replace_occured;
	main_rtio_core_outputs_collision <= 1'd0;
	main_rtio_core_outputs_collision_channel <= 1'd0;
	if ((main_rtio_core_outputs_record0_valid1 & main_rtio_core_outputs_record0_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record0_payload_channel3;
	end
	if ((main_rtio_core_outputs_record1_valid1 & main_rtio_core_outputs_record1_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record1_payload_channel3;
	end
	if ((main_rtio_core_outputs_record2_valid1 & main_rtio_core_outputs_record2_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record2_payload_channel3;
	end
	if ((main_rtio_core_outputs_record3_valid1 & main_rtio_core_outputs_record3_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record3_payload_channel3;
	end
	if ((main_rtio_core_outputs_record4_valid1 & main_rtio_core_outputs_record4_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record4_payload_channel3;
	end
	if ((main_rtio_core_outputs_record5_valid1 & main_rtio_core_outputs_record5_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record5_payload_channel3;
	end
	if ((main_rtio_core_outputs_record6_valid1 & main_rtio_core_outputs_record6_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record6_payload_channel3;
	end
	if ((main_rtio_core_outputs_record7_valid1 & main_rtio_core_outputs_record7_collision)) begin
		main_rtio_core_outputs_collision <= 1'd1;
		main_rtio_core_outputs_collision_channel <= main_rtio_core_outputs_record7_payload_channel3;
	end
	main_output_8x0_stb <= (((((((main_rtio_core_outputs_selected0 | main_rtio_core_outputs_selected1) | main_rtio_core_outputs_selected2) | main_rtio_core_outputs_selected3) | main_rtio_core_outputs_selected4) | main_rtio_core_outputs_selected5) | main_rtio_core_outputs_selected6) | main_rtio_core_outputs_selected7);
	main_output_8x0_fine_ts <= ((((((((main_rtio_core_outputs_selected0 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected1 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected2 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected3 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected4 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected5 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected6 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected7 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x0_data <= ((((((((main_rtio_core_outputs_selected0 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected1 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected2 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected3 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected4 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected5 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected6 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected7 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x1_stb <= (((((((main_rtio_core_outputs_selected8 | main_rtio_core_outputs_selected9) | main_rtio_core_outputs_selected10) | main_rtio_core_outputs_selected11) | main_rtio_core_outputs_selected12) | main_rtio_core_outputs_selected13) | main_rtio_core_outputs_selected14) | main_rtio_core_outputs_selected15);
	main_output_8x1_fine_ts <= ((((((((main_rtio_core_outputs_selected8 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected9 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected10 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected11 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected12 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected13 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected14 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected15 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x1_data <= ((((((((main_rtio_core_outputs_selected8 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected9 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected10 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected11 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected12 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected13 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected14 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected15 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x2_stb <= (((((((main_rtio_core_outputs_selected16 | main_rtio_core_outputs_selected17) | main_rtio_core_outputs_selected18) | main_rtio_core_outputs_selected19) | main_rtio_core_outputs_selected20) | main_rtio_core_outputs_selected21) | main_rtio_core_outputs_selected22) | main_rtio_core_outputs_selected23);
	main_output_8x2_fine_ts <= ((((((((main_rtio_core_outputs_selected16 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected17 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected18 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected19 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected20 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected21 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected22 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected23 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x2_data <= ((((((((main_rtio_core_outputs_selected16 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected17 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected18 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected19 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected20 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected21 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected22 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected23 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_stb <= (((((((main_rtio_core_outputs_selected24 | main_rtio_core_outputs_selected25) | main_rtio_core_outputs_selected26) | main_rtio_core_outputs_selected27) | main_rtio_core_outputs_selected28) | main_rtio_core_outputs_selected29) | main_rtio_core_outputs_selected30) | main_rtio_core_outputs_selected31);
	main_inout_8x0_inout_8x0_ointerface0_fine_ts <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_address <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x0_inout_8x0_ointerface0_data <= ((((((((main_rtio_core_outputs_selected24 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected25 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected26 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected27 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected28 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected29 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected30 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected31 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x3_stb <= (((((((main_rtio_core_outputs_selected32 | main_rtio_core_outputs_selected33) | main_rtio_core_outputs_selected34) | main_rtio_core_outputs_selected35) | main_rtio_core_outputs_selected36) | main_rtio_core_outputs_selected37) | main_rtio_core_outputs_selected38) | main_rtio_core_outputs_selected39);
	main_output_8x3_fine_ts <= ((((((((main_rtio_core_outputs_selected32 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected33 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected34 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected35 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected36 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected37 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected38 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected39 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x3_data <= ((((((((main_rtio_core_outputs_selected32 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected33 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected34 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected35 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected36 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected37 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected38 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected39 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x4_stb <= (((((((main_rtio_core_outputs_selected40 | main_rtio_core_outputs_selected41) | main_rtio_core_outputs_selected42) | main_rtio_core_outputs_selected43) | main_rtio_core_outputs_selected44) | main_rtio_core_outputs_selected45) | main_rtio_core_outputs_selected46) | main_rtio_core_outputs_selected47);
	main_output_8x4_fine_ts <= ((((((((main_rtio_core_outputs_selected40 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected41 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected42 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected43 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected44 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected45 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected46 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected47 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x4_data <= ((((((((main_rtio_core_outputs_selected40 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected41 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected42 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected43 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected44 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected45 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected46 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected47 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x5_stb <= (((((((main_rtio_core_outputs_selected48 | main_rtio_core_outputs_selected49) | main_rtio_core_outputs_selected50) | main_rtio_core_outputs_selected51) | main_rtio_core_outputs_selected52) | main_rtio_core_outputs_selected53) | main_rtio_core_outputs_selected54) | main_rtio_core_outputs_selected55);
	main_output_8x5_fine_ts <= ((((((((main_rtio_core_outputs_selected48 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected49 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected50 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected51 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected52 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected53 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected54 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected55 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x5_data <= ((((((((main_rtio_core_outputs_selected48 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected49 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected50 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected51 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected52 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected53 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected54 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected55 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_stb <= (((((((main_rtio_core_outputs_selected56 | main_rtio_core_outputs_selected57) | main_rtio_core_outputs_selected58) | main_rtio_core_outputs_selected59) | main_rtio_core_outputs_selected60) | main_rtio_core_outputs_selected61) | main_rtio_core_outputs_selected62) | main_rtio_core_outputs_selected63);
	main_inout_8x1_inout_8x1_ointerface1_fine_ts <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_address <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x1_inout_8x1_ointerface1_data <= ((((((((main_rtio_core_outputs_selected56 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected57 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected58 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected59 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected60 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected61 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected62 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected63 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x6_stb <= (((((((main_rtio_core_outputs_selected64 | main_rtio_core_outputs_selected65) | main_rtio_core_outputs_selected66) | main_rtio_core_outputs_selected67) | main_rtio_core_outputs_selected68) | main_rtio_core_outputs_selected69) | main_rtio_core_outputs_selected70) | main_rtio_core_outputs_selected71);
	main_output_8x6_fine_ts <= ((((((((main_rtio_core_outputs_selected64 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected65 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected66 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected67 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected68 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected69 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected70 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected71 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x6_data <= ((((((((main_rtio_core_outputs_selected64 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected65 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected66 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected67 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected68 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected69 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected70 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected71 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x7_stb <= (((((((main_rtio_core_outputs_selected72 | main_rtio_core_outputs_selected73) | main_rtio_core_outputs_selected74) | main_rtio_core_outputs_selected75) | main_rtio_core_outputs_selected76) | main_rtio_core_outputs_selected77) | main_rtio_core_outputs_selected78) | main_rtio_core_outputs_selected79);
	main_output_8x7_fine_ts <= ((((((((main_rtio_core_outputs_selected72 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected73 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected74 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected75 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected76 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected77 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected78 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected79 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x7_data <= ((((((((main_rtio_core_outputs_selected72 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected73 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected74 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected75 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected76 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected77 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected78 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected79 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x8_stb <= (((((((main_rtio_core_outputs_selected80 | main_rtio_core_outputs_selected81) | main_rtio_core_outputs_selected82) | main_rtio_core_outputs_selected83) | main_rtio_core_outputs_selected84) | main_rtio_core_outputs_selected85) | main_rtio_core_outputs_selected86) | main_rtio_core_outputs_selected87);
	main_output_8x8_fine_ts <= ((((((((main_rtio_core_outputs_selected80 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected81 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected82 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected83 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected84 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected85 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected86 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected87 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x8_data <= ((((((((main_rtio_core_outputs_selected80 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected81 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected82 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected83 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected84 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected85 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected86 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected87 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_stb <= (((((((main_rtio_core_outputs_selected88 | main_rtio_core_outputs_selected89) | main_rtio_core_outputs_selected90) | main_rtio_core_outputs_selected91) | main_rtio_core_outputs_selected92) | main_rtio_core_outputs_selected93) | main_rtio_core_outputs_selected94) | main_rtio_core_outputs_selected95);
	main_inout_8x2_inout_8x2_ointerface2_fine_ts <= ((((((((main_rtio_core_outputs_selected88 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected89 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected90 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected91 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected92 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected93 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected94 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected95 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_address <= ((((((((main_rtio_core_outputs_selected88 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected89 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected90 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected91 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected92 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected93 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected94 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected95 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x2_inout_8x2_ointerface2_data <= ((((((((main_rtio_core_outputs_selected88 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected89 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected90 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected91 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected92 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected93 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected94 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected95 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x9_stb <= (((((((main_rtio_core_outputs_selected96 | main_rtio_core_outputs_selected97) | main_rtio_core_outputs_selected98) | main_rtio_core_outputs_selected99) | main_rtio_core_outputs_selected100) | main_rtio_core_outputs_selected101) | main_rtio_core_outputs_selected102) | main_rtio_core_outputs_selected103);
	main_output_8x9_fine_ts <= ((((((((main_rtio_core_outputs_selected96 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected97 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected98 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected99 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected100 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected101 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected102 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected103 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x9_data <= ((((((((main_rtio_core_outputs_selected96 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected97 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected98 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected99 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected100 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected101 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected102 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected103 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x10_stb <= (((((((main_rtio_core_outputs_selected104 | main_rtio_core_outputs_selected105) | main_rtio_core_outputs_selected106) | main_rtio_core_outputs_selected107) | main_rtio_core_outputs_selected108) | main_rtio_core_outputs_selected109) | main_rtio_core_outputs_selected110) | main_rtio_core_outputs_selected111);
	main_output_8x10_fine_ts <= ((((((((main_rtio_core_outputs_selected104 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected105 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected106 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected107 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected108 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected109 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected110 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected111 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x10_data <= ((((((((main_rtio_core_outputs_selected104 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected105 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected106 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected107 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected108 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected109 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected110 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected111 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output_8x11_stb <= (((((((main_rtio_core_outputs_selected112 | main_rtio_core_outputs_selected113) | main_rtio_core_outputs_selected114) | main_rtio_core_outputs_selected115) | main_rtio_core_outputs_selected116) | main_rtio_core_outputs_selected117) | main_rtio_core_outputs_selected118) | main_rtio_core_outputs_selected119);
	main_output_8x11_fine_ts <= ((((((((main_rtio_core_outputs_selected112 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected113 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected114 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected115 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected116 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected117 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected118 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected119 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_output_8x11_data <= ((((((((main_rtio_core_outputs_selected112 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected113 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected114 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected115 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected116 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected117 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected118 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected119 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_stb <= (((((((main_rtio_core_outputs_selected120 | main_rtio_core_outputs_selected121) | main_rtio_core_outputs_selected122) | main_rtio_core_outputs_selected123) | main_rtio_core_outputs_selected124) | main_rtio_core_outputs_selected125) | main_rtio_core_outputs_selected126) | main_rtio_core_outputs_selected127);
	main_inout_8x3_inout_8x3_ointerface3_fine_ts <= ((((((((main_rtio_core_outputs_selected120 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected121 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected122 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected123 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected124 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected125 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected126 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected127 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_address <= ((((((((main_rtio_core_outputs_selected120 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected121 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected122 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected123 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected124 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected125 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected126 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected127 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x3_inout_8x3_ointerface3_data <= ((((((((main_rtio_core_outputs_selected120 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected121 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected122 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected123 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected124 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected125 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected126 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected127 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_stb <= (((((((main_rtio_core_outputs_selected128 | main_rtio_core_outputs_selected129) | main_rtio_core_outputs_selected130) | main_rtio_core_outputs_selected131) | main_rtio_core_outputs_selected132) | main_rtio_core_outputs_selected133) | main_rtio_core_outputs_selected134) | main_rtio_core_outputs_selected135);
	main_inout_8x4_inout_8x4_ointerface4_fine_ts <= ((((((((main_rtio_core_outputs_selected128 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected129 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected130 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected131 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected132 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected133 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected134 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected135 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_address <= ((((((((main_rtio_core_outputs_selected128 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected129 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected130 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected131 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected132 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected133 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected134 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected135 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x4_inout_8x4_ointerface4_data <= ((((((((main_rtio_core_outputs_selected128 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected129 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected130 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected131 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected132 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected133 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected134 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected135 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_stb <= (((((((main_rtio_core_outputs_selected136 | main_rtio_core_outputs_selected137) | main_rtio_core_outputs_selected138) | main_rtio_core_outputs_selected139) | main_rtio_core_outputs_selected140) | main_rtio_core_outputs_selected141) | main_rtio_core_outputs_selected142) | main_rtio_core_outputs_selected143);
	main_inout_8x5_inout_8x5_ointerface5_fine_ts <= ((((((((main_rtio_core_outputs_selected136 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected137 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected138 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected139 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected140 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected141 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected142 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected143 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_address <= ((((((((main_rtio_core_outputs_selected136 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected137 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected138 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected139 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected140 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected141 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected142 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected143 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x5_inout_8x5_ointerface5_data <= ((((((((main_rtio_core_outputs_selected136 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected137 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected138 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected139 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected140 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected141 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected142 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected143 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_stb <= (((((((main_rtio_core_outputs_selected144 | main_rtio_core_outputs_selected145) | main_rtio_core_outputs_selected146) | main_rtio_core_outputs_selected147) | main_rtio_core_outputs_selected148) | main_rtio_core_outputs_selected149) | main_rtio_core_outputs_selected150) | main_rtio_core_outputs_selected151);
	main_inout_8x6_inout_8x6_ointerface6_fine_ts <= ((((((((main_rtio_core_outputs_selected144 ? main_rtio_core_outputs_record0_payload_fine_ts1[2:0] : 1'd0) | (main_rtio_core_outputs_selected145 ? main_rtio_core_outputs_record1_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected146 ? main_rtio_core_outputs_record2_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected147 ? main_rtio_core_outputs_record3_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected148 ? main_rtio_core_outputs_record4_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected149 ? main_rtio_core_outputs_record5_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected150 ? main_rtio_core_outputs_record6_payload_fine_ts1[2:0] : 1'd0)) | (main_rtio_core_outputs_selected151 ? main_rtio_core_outputs_record7_payload_fine_ts1[2:0] : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_address <= ((((((((main_rtio_core_outputs_selected144 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected145 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected146 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected147 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected148 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected149 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected150 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected151 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_inout_8x6_inout_8x6_ointerface6_data <= ((((((((main_rtio_core_outputs_selected144 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected145 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected146 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected147 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected148 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected149 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected150 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected151 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output0_stb <= (((((((main_rtio_core_outputs_selected152 | main_rtio_core_outputs_selected153) | main_rtio_core_outputs_selected154) | main_rtio_core_outputs_selected155) | main_rtio_core_outputs_selected156) | main_rtio_core_outputs_selected157) | main_rtio_core_outputs_selected158) | main_rtio_core_outputs_selected159);
	main_output0_data <= ((((((((main_rtio_core_outputs_selected152 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected153 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected154 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected155 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected156 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected157 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected158 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected159 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_output1_stb <= (((((((main_rtio_core_outputs_selected160 | main_rtio_core_outputs_selected161) | main_rtio_core_outputs_selected162) | main_rtio_core_outputs_selected163) | main_rtio_core_outputs_selected164) | main_rtio_core_outputs_selected165) | main_rtio_core_outputs_selected166) | main_rtio_core_outputs_selected167);
	main_output1_data <= ((((((((main_rtio_core_outputs_selected160 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected161 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected162 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected163 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected164 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected165 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected166 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected167 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_clockgen_stb <= (((((((main_rtio_core_outputs_selected168 | main_rtio_core_outputs_selected169) | main_rtio_core_outputs_selected170) | main_rtio_core_outputs_selected171) | main_rtio_core_outputs_selected172) | main_rtio_core_outputs_selected173) | main_rtio_core_outputs_selected174) | main_rtio_core_outputs_selected175);
	main_clockgen_data <= ((((((((main_rtio_core_outputs_selected168 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected169 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected170 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected171 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected172 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected173 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected174 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected175 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster0_ointerface0_stb <= (((((((main_rtio_core_outputs_selected176 | main_rtio_core_outputs_selected177) | main_rtio_core_outputs_selected178) | main_rtio_core_outputs_selected179) | main_rtio_core_outputs_selected180) | main_rtio_core_outputs_selected181) | main_rtio_core_outputs_selected182) | main_rtio_core_outputs_selected183);
	main_spimaster0_ointerface0_address <= ((((((((main_rtio_core_outputs_selected176 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected177 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected178 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected179 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected180 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected181 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected182 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected183 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster0_ointerface0_data <= ((((((((main_rtio_core_outputs_selected176 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected177 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected178 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected179 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected180 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected181 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected182 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected183 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster1_ointerface1_stb <= (((((((main_rtio_core_outputs_selected184 | main_rtio_core_outputs_selected185) | main_rtio_core_outputs_selected186) | main_rtio_core_outputs_selected187) | main_rtio_core_outputs_selected188) | main_rtio_core_outputs_selected189) | main_rtio_core_outputs_selected190) | main_rtio_core_outputs_selected191);
	main_spimaster1_ointerface1_address <= ((((((((main_rtio_core_outputs_selected184 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected185 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected186 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected187 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected188 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected189 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected190 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected191 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster1_ointerface1_data <= ((((((((main_rtio_core_outputs_selected184 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected185 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected186 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected187 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected188 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected189 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected190 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected191 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster2_ointerface2_stb <= (((((((main_rtio_core_outputs_selected192 | main_rtio_core_outputs_selected193) | main_rtio_core_outputs_selected194) | main_rtio_core_outputs_selected195) | main_rtio_core_outputs_selected196) | main_rtio_core_outputs_selected197) | main_rtio_core_outputs_selected198) | main_rtio_core_outputs_selected199);
	main_spimaster2_ointerface2_address <= ((((((((main_rtio_core_outputs_selected192 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected193 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected194 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected195 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected196 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected197 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected198 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected199 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster2_ointerface2_data <= ((((((((main_rtio_core_outputs_selected192 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected193 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected194 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected195 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected196 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected197 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected198 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected199 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster3_ointerface3_stb <= (((((((main_rtio_core_outputs_selected200 | main_rtio_core_outputs_selected201) | main_rtio_core_outputs_selected202) | main_rtio_core_outputs_selected203) | main_rtio_core_outputs_selected204) | main_rtio_core_outputs_selected205) | main_rtio_core_outputs_selected206) | main_rtio_core_outputs_selected207);
	main_spimaster3_ointerface3_address <= ((((((((main_rtio_core_outputs_selected200 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected201 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected202 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected203 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected204 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected205 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected206 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected207 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster3_ointerface3_data <= ((((((((main_rtio_core_outputs_selected200 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected201 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected202 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected203 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected204 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected205 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected206 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected207 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_spimaster4_ointerface4_stb <= (((((((main_rtio_core_outputs_selected208 | main_rtio_core_outputs_selected209) | main_rtio_core_outputs_selected210) | main_rtio_core_outputs_selected211) | main_rtio_core_outputs_selected212) | main_rtio_core_outputs_selected213) | main_rtio_core_outputs_selected214) | main_rtio_core_outputs_selected215);
	main_spimaster4_ointerface4_address <= ((((((((main_rtio_core_outputs_selected208 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected209 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected210 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected211 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected212 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected213 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected214 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected215 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_spimaster4_ointerface4_data <= ((((((((main_rtio_core_outputs_selected208 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected209 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected210 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected211 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected212 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected213 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected214 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected215 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_ad9914_stb <= (((((((main_rtio_core_outputs_selected216 | main_rtio_core_outputs_selected217) | main_rtio_core_outputs_selected218) | main_rtio_core_outputs_selected219) | main_rtio_core_outputs_selected220) | main_rtio_core_outputs_selected221) | main_rtio_core_outputs_selected222) | main_rtio_core_outputs_selected223);
	main_ad9914_address <= ((((((((main_rtio_core_outputs_selected216 ? main_rtio_core_outputs_record0_payload_address3 : 1'd0) | (main_rtio_core_outputs_selected217 ? main_rtio_core_outputs_record1_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected218 ? main_rtio_core_outputs_record2_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected219 ? main_rtio_core_outputs_record3_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected220 ? main_rtio_core_outputs_record4_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected221 ? main_rtio_core_outputs_record5_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected222 ? main_rtio_core_outputs_record6_payload_address3 : 1'd0)) | (main_rtio_core_outputs_selected223 ? main_rtio_core_outputs_record7_payload_address3 : 1'd0));
	main_ad9914_data <= ((((((((main_rtio_core_outputs_selected216 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected217 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected218 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected219 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected220 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected221 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected222 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected223 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_stb <= (((((((main_rtio_core_outputs_selected224 | main_rtio_core_outputs_selected225) | main_rtio_core_outputs_selected226) | main_rtio_core_outputs_selected227) | main_rtio_core_outputs_selected228) | main_rtio_core_outputs_selected229) | main_rtio_core_outputs_selected230) | main_rtio_core_outputs_selected231);
	main_data <= ((((((((main_rtio_core_outputs_selected224 ? main_rtio_core_outputs_record0_payload_data3 : 1'd0) | (main_rtio_core_outputs_selected225 ? main_rtio_core_outputs_record1_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected226 ? main_rtio_core_outputs_record2_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected227 ? main_rtio_core_outputs_record3_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected228 ? main_rtio_core_outputs_record4_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected229 ? main_rtio_core_outputs_record5_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected230 ? main_rtio_core_outputs_record6_payload_data3 : 1'd0)) | (main_rtio_core_outputs_selected231 ? main_rtio_core_outputs_record7_payload_data3 : 1'd0));
	main_rtio_core_outputs_busy <= 1'd0;
	main_rtio_core_outputs_busy_channel <= 1'd0;
	main_rtio_core_outputs_stb_r0 <= (main_rtio_core_outputs_record0_valid1 & (~main_rtio_core_outputs_record0_collision));
	main_rtio_core_outputs_channel_r0 <= main_rtio_core_outputs_record0_payload_channel3;
	if ((main_rtio_core_outputs_stb_r0 & builder_sync_basiclowerer_array_muxed0)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r0;
	end
	main_rtio_core_outputs_stb_r1 <= (main_rtio_core_outputs_record1_valid1 & (~main_rtio_core_outputs_record1_collision));
	main_rtio_core_outputs_channel_r1 <= main_rtio_core_outputs_record1_payload_channel3;
	if ((main_rtio_core_outputs_stb_r1 & builder_sync_basiclowerer_array_muxed1)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r1;
	end
	main_rtio_core_outputs_stb_r2 <= (main_rtio_core_outputs_record2_valid1 & (~main_rtio_core_outputs_record2_collision));
	main_rtio_core_outputs_channel_r2 <= main_rtio_core_outputs_record2_payload_channel3;
	if ((main_rtio_core_outputs_stb_r2 & builder_sync_basiclowerer_array_muxed2)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r2;
	end
	main_rtio_core_outputs_stb_r3 <= (main_rtio_core_outputs_record3_valid1 & (~main_rtio_core_outputs_record3_collision));
	main_rtio_core_outputs_channel_r3 <= main_rtio_core_outputs_record3_payload_channel3;
	if ((main_rtio_core_outputs_stb_r3 & builder_sync_basiclowerer_array_muxed3)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r3;
	end
	main_rtio_core_outputs_stb_r4 <= (main_rtio_core_outputs_record4_valid1 & (~main_rtio_core_outputs_record4_collision));
	main_rtio_core_outputs_channel_r4 <= main_rtio_core_outputs_record4_payload_channel3;
	if ((main_rtio_core_outputs_stb_r4 & builder_sync_basiclowerer_array_muxed4)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r4;
	end
	main_rtio_core_outputs_stb_r5 <= (main_rtio_core_outputs_record5_valid1 & (~main_rtio_core_outputs_record5_collision));
	main_rtio_core_outputs_channel_r5 <= main_rtio_core_outputs_record5_payload_channel3;
	if ((main_rtio_core_outputs_stb_r5 & builder_sync_basiclowerer_array_muxed5)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r5;
	end
	main_rtio_core_outputs_stb_r6 <= (main_rtio_core_outputs_record6_valid1 & (~main_rtio_core_outputs_record6_collision));
	main_rtio_core_outputs_channel_r6 <= main_rtio_core_outputs_record6_payload_channel3;
	if ((main_rtio_core_outputs_stb_r6 & builder_sync_basiclowerer_array_muxed6)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r6;
	end
	main_rtio_core_outputs_stb_r7 <= (main_rtio_core_outputs_record7_valid1 & (~main_rtio_core_outputs_record7_collision));
	main_rtio_core_outputs_channel_r7 <= main_rtio_core_outputs_record7_payload_channel3;
	if ((main_rtio_core_outputs_stb_r7 & builder_sync_basiclowerer_array_muxed7)) begin
		main_rtio_core_outputs_busy <= 1'd1;
		main_rtio_core_outputs_busy_channel <= main_rtio_core_outputs_channel_r7;
	end
	if (({(~main_rtio_core_outputs_record0_valid0), main_rtio_core_outputs_record0_payload_channel2} == {(~main_rtio_core_outputs_record1_valid0), main_rtio_core_outputs_record1_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record0_seqn2[10] == main_rtio_core_outputs_record0_seqn2[11]) & (main_rtio_core_outputs_record1_seqn2[10] == main_rtio_core_outputs_record1_seqn2[11])) & (main_rtio_core_outputs_record0_seqn2[11] != main_rtio_core_outputs_record1_seqn2[11])) ? main_rtio_core_outputs_record0_seqn2[11] : (main_rtio_core_outputs_record0_seqn2 < main_rtio_core_outputs_record1_seqn2))) begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
		end else begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
		end
		main_rtio_core_outputs_record0_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference0;
		main_rtio_core_outputs_record1_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record0_valid0), main_rtio_core_outputs_record0_payload_channel2} < {(~main_rtio_core_outputs_record1_valid0), main_rtio_core_outputs_record1_payload_channel2})) begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
		end else begin
			main_rtio_core_outputs_record0_rec_valid <= main_rtio_core_outputs_record1_valid0;
			main_rtio_core_outputs_record0_rec_seqn <= main_rtio_core_outputs_record1_seqn2;
			main_rtio_core_outputs_record0_rec_replace_occured <= main_rtio_core_outputs_record1_replace_occured;
			main_rtio_core_outputs_record0_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_nondata_replace_occured;
			main_rtio_core_outputs_record0_rec_payload_channel <= main_rtio_core_outputs_record1_payload_channel2;
			main_rtio_core_outputs_record0_rec_payload_fine_ts <= main_rtio_core_outputs_record1_payload_fine_ts0;
			main_rtio_core_outputs_record0_rec_payload_address <= main_rtio_core_outputs_record1_payload_address2;
			main_rtio_core_outputs_record0_rec_payload_data <= main_rtio_core_outputs_record1_payload_data2;
			main_rtio_core_outputs_record1_rec_valid <= main_rtio_core_outputs_record0_valid0;
			main_rtio_core_outputs_record1_rec_seqn <= main_rtio_core_outputs_record0_seqn2;
			main_rtio_core_outputs_record1_rec_replace_occured <= main_rtio_core_outputs_record0_replace_occured;
			main_rtio_core_outputs_record1_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_nondata_replace_occured;
			main_rtio_core_outputs_record1_rec_payload_channel <= main_rtio_core_outputs_record0_payload_channel2;
			main_rtio_core_outputs_record1_rec_payload_fine_ts <= main_rtio_core_outputs_record0_payload_fine_ts0;
			main_rtio_core_outputs_record1_rec_payload_address <= main_rtio_core_outputs_record0_payload_address2;
			main_rtio_core_outputs_record1_rec_payload_data <= main_rtio_core_outputs_record0_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record2_valid0), main_rtio_core_outputs_record2_payload_channel2} == {(~main_rtio_core_outputs_record3_valid0), main_rtio_core_outputs_record3_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record2_seqn2[10] == main_rtio_core_outputs_record2_seqn2[11]) & (main_rtio_core_outputs_record3_seqn2[10] == main_rtio_core_outputs_record3_seqn2[11])) & (main_rtio_core_outputs_record2_seqn2[11] != main_rtio_core_outputs_record3_seqn2[11])) ? main_rtio_core_outputs_record2_seqn2[11] : (main_rtio_core_outputs_record2_seqn2 < main_rtio_core_outputs_record3_seqn2))) begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
		end else begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
		end
		main_rtio_core_outputs_record2_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference1;
		main_rtio_core_outputs_record3_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record2_valid0), main_rtio_core_outputs_record2_payload_channel2} < {(~main_rtio_core_outputs_record3_valid0), main_rtio_core_outputs_record3_payload_channel2})) begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
		end else begin
			main_rtio_core_outputs_record2_rec_valid <= main_rtio_core_outputs_record3_valid0;
			main_rtio_core_outputs_record2_rec_seqn <= main_rtio_core_outputs_record3_seqn2;
			main_rtio_core_outputs_record2_rec_replace_occured <= main_rtio_core_outputs_record3_replace_occured;
			main_rtio_core_outputs_record2_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_nondata_replace_occured;
			main_rtio_core_outputs_record2_rec_payload_channel <= main_rtio_core_outputs_record3_payload_channel2;
			main_rtio_core_outputs_record2_rec_payload_fine_ts <= main_rtio_core_outputs_record3_payload_fine_ts0;
			main_rtio_core_outputs_record2_rec_payload_address <= main_rtio_core_outputs_record3_payload_address2;
			main_rtio_core_outputs_record2_rec_payload_data <= main_rtio_core_outputs_record3_payload_data2;
			main_rtio_core_outputs_record3_rec_valid <= main_rtio_core_outputs_record2_valid0;
			main_rtio_core_outputs_record3_rec_seqn <= main_rtio_core_outputs_record2_seqn2;
			main_rtio_core_outputs_record3_rec_replace_occured <= main_rtio_core_outputs_record2_replace_occured;
			main_rtio_core_outputs_record3_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_nondata_replace_occured;
			main_rtio_core_outputs_record3_rec_payload_channel <= main_rtio_core_outputs_record2_payload_channel2;
			main_rtio_core_outputs_record3_rec_payload_fine_ts <= main_rtio_core_outputs_record2_payload_fine_ts0;
			main_rtio_core_outputs_record3_rec_payload_address <= main_rtio_core_outputs_record2_payload_address2;
			main_rtio_core_outputs_record3_rec_payload_data <= main_rtio_core_outputs_record2_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record4_valid0), main_rtio_core_outputs_record4_payload_channel2} == {(~main_rtio_core_outputs_record5_valid0), main_rtio_core_outputs_record5_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record4_seqn2[10] == main_rtio_core_outputs_record4_seqn2[11]) & (main_rtio_core_outputs_record5_seqn2[10] == main_rtio_core_outputs_record5_seqn2[11])) & (main_rtio_core_outputs_record4_seqn2[11] != main_rtio_core_outputs_record5_seqn2[11])) ? main_rtio_core_outputs_record4_seqn2[11] : (main_rtio_core_outputs_record4_seqn2 < main_rtio_core_outputs_record5_seqn2))) begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
		end else begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
		end
		main_rtio_core_outputs_record4_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference2;
		main_rtio_core_outputs_record5_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record4_valid0), main_rtio_core_outputs_record4_payload_channel2} < {(~main_rtio_core_outputs_record5_valid0), main_rtio_core_outputs_record5_payload_channel2})) begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
		end else begin
			main_rtio_core_outputs_record4_rec_valid <= main_rtio_core_outputs_record5_valid0;
			main_rtio_core_outputs_record4_rec_seqn <= main_rtio_core_outputs_record5_seqn2;
			main_rtio_core_outputs_record4_rec_replace_occured <= main_rtio_core_outputs_record5_replace_occured;
			main_rtio_core_outputs_record4_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_nondata_replace_occured;
			main_rtio_core_outputs_record4_rec_payload_channel <= main_rtio_core_outputs_record5_payload_channel2;
			main_rtio_core_outputs_record4_rec_payload_fine_ts <= main_rtio_core_outputs_record5_payload_fine_ts0;
			main_rtio_core_outputs_record4_rec_payload_address <= main_rtio_core_outputs_record5_payload_address2;
			main_rtio_core_outputs_record4_rec_payload_data <= main_rtio_core_outputs_record5_payload_data2;
			main_rtio_core_outputs_record5_rec_valid <= main_rtio_core_outputs_record4_valid0;
			main_rtio_core_outputs_record5_rec_seqn <= main_rtio_core_outputs_record4_seqn2;
			main_rtio_core_outputs_record5_rec_replace_occured <= main_rtio_core_outputs_record4_replace_occured;
			main_rtio_core_outputs_record5_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_nondata_replace_occured;
			main_rtio_core_outputs_record5_rec_payload_channel <= main_rtio_core_outputs_record4_payload_channel2;
			main_rtio_core_outputs_record5_rec_payload_fine_ts <= main_rtio_core_outputs_record4_payload_fine_ts0;
			main_rtio_core_outputs_record5_rec_payload_address <= main_rtio_core_outputs_record4_payload_address2;
			main_rtio_core_outputs_record5_rec_payload_data <= main_rtio_core_outputs_record4_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record6_valid0), main_rtio_core_outputs_record6_payload_channel2} == {(~main_rtio_core_outputs_record7_valid0), main_rtio_core_outputs_record7_payload_channel2})) begin
		if (((((main_rtio_core_outputs_record6_seqn2[10] == main_rtio_core_outputs_record6_seqn2[11]) & (main_rtio_core_outputs_record7_seqn2[10] == main_rtio_core_outputs_record7_seqn2[11])) & (main_rtio_core_outputs_record6_seqn2[11] != main_rtio_core_outputs_record7_seqn2[11])) ? main_rtio_core_outputs_record6_seqn2[11] : (main_rtio_core_outputs_record6_seqn2 < main_rtio_core_outputs_record7_seqn2))) begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
		end else begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
		end
		main_rtio_core_outputs_record6_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference3;
		main_rtio_core_outputs_record7_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record6_valid0), main_rtio_core_outputs_record6_payload_channel2} < {(~main_rtio_core_outputs_record7_valid0), main_rtio_core_outputs_record7_payload_channel2})) begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
		end else begin
			main_rtio_core_outputs_record6_rec_valid <= main_rtio_core_outputs_record7_valid0;
			main_rtio_core_outputs_record6_rec_seqn <= main_rtio_core_outputs_record7_seqn2;
			main_rtio_core_outputs_record6_rec_replace_occured <= main_rtio_core_outputs_record7_replace_occured;
			main_rtio_core_outputs_record6_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_nondata_replace_occured;
			main_rtio_core_outputs_record6_rec_payload_channel <= main_rtio_core_outputs_record7_payload_channel2;
			main_rtio_core_outputs_record6_rec_payload_fine_ts <= main_rtio_core_outputs_record7_payload_fine_ts0;
			main_rtio_core_outputs_record6_rec_payload_address <= main_rtio_core_outputs_record7_payload_address2;
			main_rtio_core_outputs_record6_rec_payload_data <= main_rtio_core_outputs_record7_payload_data2;
			main_rtio_core_outputs_record7_rec_valid <= main_rtio_core_outputs_record6_valid0;
			main_rtio_core_outputs_record7_rec_seqn <= main_rtio_core_outputs_record6_seqn2;
			main_rtio_core_outputs_record7_rec_replace_occured <= main_rtio_core_outputs_record6_replace_occured;
			main_rtio_core_outputs_record7_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_nondata_replace_occured;
			main_rtio_core_outputs_record7_rec_payload_channel <= main_rtio_core_outputs_record6_payload_channel2;
			main_rtio_core_outputs_record7_rec_payload_fine_ts <= main_rtio_core_outputs_record6_payload_fine_ts0;
			main_rtio_core_outputs_record7_rec_payload_address <= main_rtio_core_outputs_record6_payload_address2;
			main_rtio_core_outputs_record7_rec_payload_data <= main_rtio_core_outputs_record6_payload_data2;
		end
	end
	if (({(~main_rtio_core_outputs_record0_rec_valid), main_rtio_core_outputs_record0_rec_payload_channel} == {(~main_rtio_core_outputs_record2_rec_valid), main_rtio_core_outputs_record2_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record0_rec_seqn[10] == main_rtio_core_outputs_record0_rec_seqn[11]) & (main_rtio_core_outputs_record2_rec_seqn[10] == main_rtio_core_outputs_record2_rec_seqn[11])) & (main_rtio_core_outputs_record0_rec_seqn[11] != main_rtio_core_outputs_record2_rec_seqn[11])) ? main_rtio_core_outputs_record0_rec_seqn[11] : (main_rtio_core_outputs_record0_rec_seqn < main_rtio_core_outputs_record2_rec_seqn))) begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
		end
		main_rtio_core_outputs_record8_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference4;
		main_rtio_core_outputs_record10_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record0_rec_valid), main_rtio_core_outputs_record0_rec_payload_channel} < {(~main_rtio_core_outputs_record2_rec_valid), main_rtio_core_outputs_record2_rec_payload_channel})) begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record8_rec_valid <= main_rtio_core_outputs_record2_rec_valid;
			main_rtio_core_outputs_record8_rec_seqn <= main_rtio_core_outputs_record2_rec_seqn;
			main_rtio_core_outputs_record8_rec_replace_occured <= main_rtio_core_outputs_record2_rec_replace_occured;
			main_rtio_core_outputs_record8_rec_nondata_replace_occured <= main_rtio_core_outputs_record2_rec_nondata_replace_occured;
			main_rtio_core_outputs_record8_rec_payload_channel <= main_rtio_core_outputs_record2_rec_payload_channel;
			main_rtio_core_outputs_record8_rec_payload_fine_ts <= main_rtio_core_outputs_record2_rec_payload_fine_ts;
			main_rtio_core_outputs_record8_rec_payload_address <= main_rtio_core_outputs_record2_rec_payload_address;
			main_rtio_core_outputs_record8_rec_payload_data <= main_rtio_core_outputs_record2_rec_payload_data;
			main_rtio_core_outputs_record10_rec_valid <= main_rtio_core_outputs_record0_rec_valid;
			main_rtio_core_outputs_record10_rec_seqn <= main_rtio_core_outputs_record0_rec_seqn;
			main_rtio_core_outputs_record10_rec_replace_occured <= main_rtio_core_outputs_record0_rec_replace_occured;
			main_rtio_core_outputs_record10_rec_nondata_replace_occured <= main_rtio_core_outputs_record0_rec_nondata_replace_occured;
			main_rtio_core_outputs_record10_rec_payload_channel <= main_rtio_core_outputs_record0_rec_payload_channel;
			main_rtio_core_outputs_record10_rec_payload_fine_ts <= main_rtio_core_outputs_record0_rec_payload_fine_ts;
			main_rtio_core_outputs_record10_rec_payload_address <= main_rtio_core_outputs_record0_rec_payload_address;
			main_rtio_core_outputs_record10_rec_payload_data <= main_rtio_core_outputs_record0_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record1_rec_valid), main_rtio_core_outputs_record1_rec_payload_channel} == {(~main_rtio_core_outputs_record3_rec_valid), main_rtio_core_outputs_record3_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record1_rec_seqn[10] == main_rtio_core_outputs_record1_rec_seqn[11]) & (main_rtio_core_outputs_record3_rec_seqn[10] == main_rtio_core_outputs_record3_rec_seqn[11])) & (main_rtio_core_outputs_record1_rec_seqn[11] != main_rtio_core_outputs_record3_rec_seqn[11])) ? main_rtio_core_outputs_record1_rec_seqn[11] : (main_rtio_core_outputs_record1_rec_seqn < main_rtio_core_outputs_record3_rec_seqn))) begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
		end
		main_rtio_core_outputs_record9_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference5;
		main_rtio_core_outputs_record11_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record1_rec_valid), main_rtio_core_outputs_record1_rec_payload_channel} < {(~main_rtio_core_outputs_record3_rec_valid), main_rtio_core_outputs_record3_rec_payload_channel})) begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record9_rec_valid <= main_rtio_core_outputs_record3_rec_valid;
			main_rtio_core_outputs_record9_rec_seqn <= main_rtio_core_outputs_record3_rec_seqn;
			main_rtio_core_outputs_record9_rec_replace_occured <= main_rtio_core_outputs_record3_rec_replace_occured;
			main_rtio_core_outputs_record9_rec_nondata_replace_occured <= main_rtio_core_outputs_record3_rec_nondata_replace_occured;
			main_rtio_core_outputs_record9_rec_payload_channel <= main_rtio_core_outputs_record3_rec_payload_channel;
			main_rtio_core_outputs_record9_rec_payload_fine_ts <= main_rtio_core_outputs_record3_rec_payload_fine_ts;
			main_rtio_core_outputs_record9_rec_payload_address <= main_rtio_core_outputs_record3_rec_payload_address;
			main_rtio_core_outputs_record9_rec_payload_data <= main_rtio_core_outputs_record3_rec_payload_data;
			main_rtio_core_outputs_record11_rec_valid <= main_rtio_core_outputs_record1_rec_valid;
			main_rtio_core_outputs_record11_rec_seqn <= main_rtio_core_outputs_record1_rec_seqn;
			main_rtio_core_outputs_record11_rec_replace_occured <= main_rtio_core_outputs_record1_rec_replace_occured;
			main_rtio_core_outputs_record11_rec_nondata_replace_occured <= main_rtio_core_outputs_record1_rec_nondata_replace_occured;
			main_rtio_core_outputs_record11_rec_payload_channel <= main_rtio_core_outputs_record1_rec_payload_channel;
			main_rtio_core_outputs_record11_rec_payload_fine_ts <= main_rtio_core_outputs_record1_rec_payload_fine_ts;
			main_rtio_core_outputs_record11_rec_payload_address <= main_rtio_core_outputs_record1_rec_payload_address;
			main_rtio_core_outputs_record11_rec_payload_data <= main_rtio_core_outputs_record1_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record4_rec_valid), main_rtio_core_outputs_record4_rec_payload_channel} == {(~main_rtio_core_outputs_record6_rec_valid), main_rtio_core_outputs_record6_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record4_rec_seqn[10] == main_rtio_core_outputs_record4_rec_seqn[11]) & (main_rtio_core_outputs_record6_rec_seqn[10] == main_rtio_core_outputs_record6_rec_seqn[11])) & (main_rtio_core_outputs_record4_rec_seqn[11] != main_rtio_core_outputs_record6_rec_seqn[11])) ? main_rtio_core_outputs_record4_rec_seqn[11] : (main_rtio_core_outputs_record4_rec_seqn < main_rtio_core_outputs_record6_rec_seqn))) begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
		end
		main_rtio_core_outputs_record12_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference6;
		main_rtio_core_outputs_record14_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record4_rec_valid), main_rtio_core_outputs_record4_rec_payload_channel} < {(~main_rtio_core_outputs_record6_rec_valid), main_rtio_core_outputs_record6_rec_payload_channel})) begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record12_rec_valid <= main_rtio_core_outputs_record6_rec_valid;
			main_rtio_core_outputs_record12_rec_seqn <= main_rtio_core_outputs_record6_rec_seqn;
			main_rtio_core_outputs_record12_rec_replace_occured <= main_rtio_core_outputs_record6_rec_replace_occured;
			main_rtio_core_outputs_record12_rec_nondata_replace_occured <= main_rtio_core_outputs_record6_rec_nondata_replace_occured;
			main_rtio_core_outputs_record12_rec_payload_channel <= main_rtio_core_outputs_record6_rec_payload_channel;
			main_rtio_core_outputs_record12_rec_payload_fine_ts <= main_rtio_core_outputs_record6_rec_payload_fine_ts;
			main_rtio_core_outputs_record12_rec_payload_address <= main_rtio_core_outputs_record6_rec_payload_address;
			main_rtio_core_outputs_record12_rec_payload_data <= main_rtio_core_outputs_record6_rec_payload_data;
			main_rtio_core_outputs_record14_rec_valid <= main_rtio_core_outputs_record4_rec_valid;
			main_rtio_core_outputs_record14_rec_seqn <= main_rtio_core_outputs_record4_rec_seqn;
			main_rtio_core_outputs_record14_rec_replace_occured <= main_rtio_core_outputs_record4_rec_replace_occured;
			main_rtio_core_outputs_record14_rec_nondata_replace_occured <= main_rtio_core_outputs_record4_rec_nondata_replace_occured;
			main_rtio_core_outputs_record14_rec_payload_channel <= main_rtio_core_outputs_record4_rec_payload_channel;
			main_rtio_core_outputs_record14_rec_payload_fine_ts <= main_rtio_core_outputs_record4_rec_payload_fine_ts;
			main_rtio_core_outputs_record14_rec_payload_address <= main_rtio_core_outputs_record4_rec_payload_address;
			main_rtio_core_outputs_record14_rec_payload_data <= main_rtio_core_outputs_record4_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record5_rec_valid), main_rtio_core_outputs_record5_rec_payload_channel} == {(~main_rtio_core_outputs_record7_rec_valid), main_rtio_core_outputs_record7_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record5_rec_seqn[10] == main_rtio_core_outputs_record5_rec_seqn[11]) & (main_rtio_core_outputs_record7_rec_seqn[10] == main_rtio_core_outputs_record7_rec_seqn[11])) & (main_rtio_core_outputs_record5_rec_seqn[11] != main_rtio_core_outputs_record7_rec_seqn[11])) ? main_rtio_core_outputs_record5_rec_seqn[11] : (main_rtio_core_outputs_record5_rec_seqn < main_rtio_core_outputs_record7_rec_seqn))) begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
		end
		main_rtio_core_outputs_record13_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference7;
		main_rtio_core_outputs_record15_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record5_rec_valid), main_rtio_core_outputs_record5_rec_payload_channel} < {(~main_rtio_core_outputs_record7_rec_valid), main_rtio_core_outputs_record7_rec_payload_channel})) begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record13_rec_valid <= main_rtio_core_outputs_record7_rec_valid;
			main_rtio_core_outputs_record13_rec_seqn <= main_rtio_core_outputs_record7_rec_seqn;
			main_rtio_core_outputs_record13_rec_replace_occured <= main_rtio_core_outputs_record7_rec_replace_occured;
			main_rtio_core_outputs_record13_rec_nondata_replace_occured <= main_rtio_core_outputs_record7_rec_nondata_replace_occured;
			main_rtio_core_outputs_record13_rec_payload_channel <= main_rtio_core_outputs_record7_rec_payload_channel;
			main_rtio_core_outputs_record13_rec_payload_fine_ts <= main_rtio_core_outputs_record7_rec_payload_fine_ts;
			main_rtio_core_outputs_record13_rec_payload_address <= main_rtio_core_outputs_record7_rec_payload_address;
			main_rtio_core_outputs_record13_rec_payload_data <= main_rtio_core_outputs_record7_rec_payload_data;
			main_rtio_core_outputs_record15_rec_valid <= main_rtio_core_outputs_record5_rec_valid;
			main_rtio_core_outputs_record15_rec_seqn <= main_rtio_core_outputs_record5_rec_seqn;
			main_rtio_core_outputs_record15_rec_replace_occured <= main_rtio_core_outputs_record5_rec_replace_occured;
			main_rtio_core_outputs_record15_rec_nondata_replace_occured <= main_rtio_core_outputs_record5_rec_nondata_replace_occured;
			main_rtio_core_outputs_record15_rec_payload_channel <= main_rtio_core_outputs_record5_rec_payload_channel;
			main_rtio_core_outputs_record15_rec_payload_fine_ts <= main_rtio_core_outputs_record5_rec_payload_fine_ts;
			main_rtio_core_outputs_record15_rec_payload_address <= main_rtio_core_outputs_record5_rec_payload_address;
			main_rtio_core_outputs_record15_rec_payload_data <= main_rtio_core_outputs_record5_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record9_rec_valid), main_rtio_core_outputs_record9_rec_payload_channel} == {(~main_rtio_core_outputs_record10_rec_valid), main_rtio_core_outputs_record10_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record9_rec_seqn[10] == main_rtio_core_outputs_record9_rec_seqn[11]) & (main_rtio_core_outputs_record10_rec_seqn[10] == main_rtio_core_outputs_record10_rec_seqn[11])) & (main_rtio_core_outputs_record9_rec_seqn[11] != main_rtio_core_outputs_record10_rec_seqn[11])) ? main_rtio_core_outputs_record9_rec_seqn[11] : (main_rtio_core_outputs_record9_rec_seqn < main_rtio_core_outputs_record10_rec_seqn))) begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
		end
		main_rtio_core_outputs_record17_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference8;
		main_rtio_core_outputs_record18_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record9_rec_valid), main_rtio_core_outputs_record9_rec_payload_channel} < {(~main_rtio_core_outputs_record10_rec_valid), main_rtio_core_outputs_record10_rec_payload_channel})) begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record17_rec_valid <= main_rtio_core_outputs_record10_rec_valid;
			main_rtio_core_outputs_record17_rec_seqn <= main_rtio_core_outputs_record10_rec_seqn;
			main_rtio_core_outputs_record17_rec_replace_occured <= main_rtio_core_outputs_record10_rec_replace_occured;
			main_rtio_core_outputs_record17_rec_nondata_replace_occured <= main_rtio_core_outputs_record10_rec_nondata_replace_occured;
			main_rtio_core_outputs_record17_rec_payload_channel <= main_rtio_core_outputs_record10_rec_payload_channel;
			main_rtio_core_outputs_record17_rec_payload_fine_ts <= main_rtio_core_outputs_record10_rec_payload_fine_ts;
			main_rtio_core_outputs_record17_rec_payload_address <= main_rtio_core_outputs_record10_rec_payload_address;
			main_rtio_core_outputs_record17_rec_payload_data <= main_rtio_core_outputs_record10_rec_payload_data;
			main_rtio_core_outputs_record18_rec_valid <= main_rtio_core_outputs_record9_rec_valid;
			main_rtio_core_outputs_record18_rec_seqn <= main_rtio_core_outputs_record9_rec_seqn;
			main_rtio_core_outputs_record18_rec_replace_occured <= main_rtio_core_outputs_record9_rec_replace_occured;
			main_rtio_core_outputs_record18_rec_nondata_replace_occured <= main_rtio_core_outputs_record9_rec_nondata_replace_occured;
			main_rtio_core_outputs_record18_rec_payload_channel <= main_rtio_core_outputs_record9_rec_payload_channel;
			main_rtio_core_outputs_record18_rec_payload_fine_ts <= main_rtio_core_outputs_record9_rec_payload_fine_ts;
			main_rtio_core_outputs_record18_rec_payload_address <= main_rtio_core_outputs_record9_rec_payload_address;
			main_rtio_core_outputs_record18_rec_payload_data <= main_rtio_core_outputs_record9_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record13_rec_valid), main_rtio_core_outputs_record13_rec_payload_channel} == {(~main_rtio_core_outputs_record14_rec_valid), main_rtio_core_outputs_record14_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record13_rec_seqn[10] == main_rtio_core_outputs_record13_rec_seqn[11]) & (main_rtio_core_outputs_record14_rec_seqn[10] == main_rtio_core_outputs_record14_rec_seqn[11])) & (main_rtio_core_outputs_record13_rec_seqn[11] != main_rtio_core_outputs_record14_rec_seqn[11])) ? main_rtio_core_outputs_record13_rec_seqn[11] : (main_rtio_core_outputs_record13_rec_seqn < main_rtio_core_outputs_record14_rec_seqn))) begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
		end
		main_rtio_core_outputs_record21_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference9;
		main_rtio_core_outputs_record22_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record13_rec_valid), main_rtio_core_outputs_record13_rec_payload_channel} < {(~main_rtio_core_outputs_record14_rec_valid), main_rtio_core_outputs_record14_rec_payload_channel})) begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record21_rec_valid <= main_rtio_core_outputs_record14_rec_valid;
			main_rtio_core_outputs_record21_rec_seqn <= main_rtio_core_outputs_record14_rec_seqn;
			main_rtio_core_outputs_record21_rec_replace_occured <= main_rtio_core_outputs_record14_rec_replace_occured;
			main_rtio_core_outputs_record21_rec_nondata_replace_occured <= main_rtio_core_outputs_record14_rec_nondata_replace_occured;
			main_rtio_core_outputs_record21_rec_payload_channel <= main_rtio_core_outputs_record14_rec_payload_channel;
			main_rtio_core_outputs_record21_rec_payload_fine_ts <= main_rtio_core_outputs_record14_rec_payload_fine_ts;
			main_rtio_core_outputs_record21_rec_payload_address <= main_rtio_core_outputs_record14_rec_payload_address;
			main_rtio_core_outputs_record21_rec_payload_data <= main_rtio_core_outputs_record14_rec_payload_data;
			main_rtio_core_outputs_record22_rec_valid <= main_rtio_core_outputs_record13_rec_valid;
			main_rtio_core_outputs_record22_rec_seqn <= main_rtio_core_outputs_record13_rec_seqn;
			main_rtio_core_outputs_record22_rec_replace_occured <= main_rtio_core_outputs_record13_rec_replace_occured;
			main_rtio_core_outputs_record22_rec_nondata_replace_occured <= main_rtio_core_outputs_record13_rec_nondata_replace_occured;
			main_rtio_core_outputs_record22_rec_payload_channel <= main_rtio_core_outputs_record13_rec_payload_channel;
			main_rtio_core_outputs_record22_rec_payload_fine_ts <= main_rtio_core_outputs_record13_rec_payload_fine_ts;
			main_rtio_core_outputs_record22_rec_payload_address <= main_rtio_core_outputs_record13_rec_payload_address;
			main_rtio_core_outputs_record22_rec_payload_data <= main_rtio_core_outputs_record13_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record16_rec_valid <= main_rtio_core_outputs_record8_rec_valid;
	main_rtio_core_outputs_record16_rec_seqn <= main_rtio_core_outputs_record8_rec_seqn;
	main_rtio_core_outputs_record16_rec_replace_occured <= main_rtio_core_outputs_record8_rec_replace_occured;
	main_rtio_core_outputs_record16_rec_nondata_replace_occured <= main_rtio_core_outputs_record8_rec_nondata_replace_occured;
	main_rtio_core_outputs_record16_rec_payload_channel <= main_rtio_core_outputs_record8_rec_payload_channel;
	main_rtio_core_outputs_record16_rec_payload_fine_ts <= main_rtio_core_outputs_record8_rec_payload_fine_ts;
	main_rtio_core_outputs_record16_rec_payload_address <= main_rtio_core_outputs_record8_rec_payload_address;
	main_rtio_core_outputs_record16_rec_payload_data <= main_rtio_core_outputs_record8_rec_payload_data;
	main_rtio_core_outputs_record19_rec_valid <= main_rtio_core_outputs_record11_rec_valid;
	main_rtio_core_outputs_record19_rec_seqn <= main_rtio_core_outputs_record11_rec_seqn;
	main_rtio_core_outputs_record19_rec_replace_occured <= main_rtio_core_outputs_record11_rec_replace_occured;
	main_rtio_core_outputs_record19_rec_nondata_replace_occured <= main_rtio_core_outputs_record11_rec_nondata_replace_occured;
	main_rtio_core_outputs_record19_rec_payload_channel <= main_rtio_core_outputs_record11_rec_payload_channel;
	main_rtio_core_outputs_record19_rec_payload_fine_ts <= main_rtio_core_outputs_record11_rec_payload_fine_ts;
	main_rtio_core_outputs_record19_rec_payload_address <= main_rtio_core_outputs_record11_rec_payload_address;
	main_rtio_core_outputs_record19_rec_payload_data <= main_rtio_core_outputs_record11_rec_payload_data;
	main_rtio_core_outputs_record20_rec_valid <= main_rtio_core_outputs_record12_rec_valid;
	main_rtio_core_outputs_record20_rec_seqn <= main_rtio_core_outputs_record12_rec_seqn;
	main_rtio_core_outputs_record20_rec_replace_occured <= main_rtio_core_outputs_record12_rec_replace_occured;
	main_rtio_core_outputs_record20_rec_nondata_replace_occured <= main_rtio_core_outputs_record12_rec_nondata_replace_occured;
	main_rtio_core_outputs_record20_rec_payload_channel <= main_rtio_core_outputs_record12_rec_payload_channel;
	main_rtio_core_outputs_record20_rec_payload_fine_ts <= main_rtio_core_outputs_record12_rec_payload_fine_ts;
	main_rtio_core_outputs_record20_rec_payload_address <= main_rtio_core_outputs_record12_rec_payload_address;
	main_rtio_core_outputs_record20_rec_payload_data <= main_rtio_core_outputs_record12_rec_payload_data;
	main_rtio_core_outputs_record23_rec_valid <= main_rtio_core_outputs_record15_rec_valid;
	main_rtio_core_outputs_record23_rec_seqn <= main_rtio_core_outputs_record15_rec_seqn;
	main_rtio_core_outputs_record23_rec_replace_occured <= main_rtio_core_outputs_record15_rec_replace_occured;
	main_rtio_core_outputs_record23_rec_nondata_replace_occured <= main_rtio_core_outputs_record15_rec_nondata_replace_occured;
	main_rtio_core_outputs_record23_rec_payload_channel <= main_rtio_core_outputs_record15_rec_payload_channel;
	main_rtio_core_outputs_record23_rec_payload_fine_ts <= main_rtio_core_outputs_record15_rec_payload_fine_ts;
	main_rtio_core_outputs_record23_rec_payload_address <= main_rtio_core_outputs_record15_rec_payload_address;
	main_rtio_core_outputs_record23_rec_payload_data <= main_rtio_core_outputs_record15_rec_payload_data;
	if (({(~main_rtio_core_outputs_record16_rec_valid), main_rtio_core_outputs_record16_rec_payload_channel} == {(~main_rtio_core_outputs_record20_rec_valid), main_rtio_core_outputs_record20_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record16_rec_seqn[10] == main_rtio_core_outputs_record16_rec_seqn[11]) & (main_rtio_core_outputs_record20_rec_seqn[10] == main_rtio_core_outputs_record20_rec_seqn[11])) & (main_rtio_core_outputs_record16_rec_seqn[11] != main_rtio_core_outputs_record20_rec_seqn[11])) ? main_rtio_core_outputs_record16_rec_seqn[11] : (main_rtio_core_outputs_record16_rec_seqn < main_rtio_core_outputs_record20_rec_seqn))) begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
		end
		main_rtio_core_outputs_record24_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference10;
		main_rtio_core_outputs_record28_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record16_rec_valid), main_rtio_core_outputs_record16_rec_payload_channel} < {(~main_rtio_core_outputs_record20_rec_valid), main_rtio_core_outputs_record20_rec_payload_channel})) begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record24_rec_valid <= main_rtio_core_outputs_record20_rec_valid;
			main_rtio_core_outputs_record24_rec_seqn <= main_rtio_core_outputs_record20_rec_seqn;
			main_rtio_core_outputs_record24_rec_replace_occured <= main_rtio_core_outputs_record20_rec_replace_occured;
			main_rtio_core_outputs_record24_rec_nondata_replace_occured <= main_rtio_core_outputs_record20_rec_nondata_replace_occured;
			main_rtio_core_outputs_record24_rec_payload_channel <= main_rtio_core_outputs_record20_rec_payload_channel;
			main_rtio_core_outputs_record24_rec_payload_fine_ts <= main_rtio_core_outputs_record20_rec_payload_fine_ts;
			main_rtio_core_outputs_record24_rec_payload_address <= main_rtio_core_outputs_record20_rec_payload_address;
			main_rtio_core_outputs_record24_rec_payload_data <= main_rtio_core_outputs_record20_rec_payload_data;
			main_rtio_core_outputs_record28_rec_valid <= main_rtio_core_outputs_record16_rec_valid;
			main_rtio_core_outputs_record28_rec_seqn <= main_rtio_core_outputs_record16_rec_seqn;
			main_rtio_core_outputs_record28_rec_replace_occured <= main_rtio_core_outputs_record16_rec_replace_occured;
			main_rtio_core_outputs_record28_rec_nondata_replace_occured <= main_rtio_core_outputs_record16_rec_nondata_replace_occured;
			main_rtio_core_outputs_record28_rec_payload_channel <= main_rtio_core_outputs_record16_rec_payload_channel;
			main_rtio_core_outputs_record28_rec_payload_fine_ts <= main_rtio_core_outputs_record16_rec_payload_fine_ts;
			main_rtio_core_outputs_record28_rec_payload_address <= main_rtio_core_outputs_record16_rec_payload_address;
			main_rtio_core_outputs_record28_rec_payload_data <= main_rtio_core_outputs_record16_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record17_rec_valid), main_rtio_core_outputs_record17_rec_payload_channel} == {(~main_rtio_core_outputs_record21_rec_valid), main_rtio_core_outputs_record21_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record17_rec_seqn[10] == main_rtio_core_outputs_record17_rec_seqn[11]) & (main_rtio_core_outputs_record21_rec_seqn[10] == main_rtio_core_outputs_record21_rec_seqn[11])) & (main_rtio_core_outputs_record17_rec_seqn[11] != main_rtio_core_outputs_record21_rec_seqn[11])) ? main_rtio_core_outputs_record17_rec_seqn[11] : (main_rtio_core_outputs_record17_rec_seqn < main_rtio_core_outputs_record21_rec_seqn))) begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
		end
		main_rtio_core_outputs_record25_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference11;
		main_rtio_core_outputs_record29_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record17_rec_valid), main_rtio_core_outputs_record17_rec_payload_channel} < {(~main_rtio_core_outputs_record21_rec_valid), main_rtio_core_outputs_record21_rec_payload_channel})) begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record25_rec_valid <= main_rtio_core_outputs_record21_rec_valid;
			main_rtio_core_outputs_record25_rec_seqn <= main_rtio_core_outputs_record21_rec_seqn;
			main_rtio_core_outputs_record25_rec_replace_occured <= main_rtio_core_outputs_record21_rec_replace_occured;
			main_rtio_core_outputs_record25_rec_nondata_replace_occured <= main_rtio_core_outputs_record21_rec_nondata_replace_occured;
			main_rtio_core_outputs_record25_rec_payload_channel <= main_rtio_core_outputs_record21_rec_payload_channel;
			main_rtio_core_outputs_record25_rec_payload_fine_ts <= main_rtio_core_outputs_record21_rec_payload_fine_ts;
			main_rtio_core_outputs_record25_rec_payload_address <= main_rtio_core_outputs_record21_rec_payload_address;
			main_rtio_core_outputs_record25_rec_payload_data <= main_rtio_core_outputs_record21_rec_payload_data;
			main_rtio_core_outputs_record29_rec_valid <= main_rtio_core_outputs_record17_rec_valid;
			main_rtio_core_outputs_record29_rec_seqn <= main_rtio_core_outputs_record17_rec_seqn;
			main_rtio_core_outputs_record29_rec_replace_occured <= main_rtio_core_outputs_record17_rec_replace_occured;
			main_rtio_core_outputs_record29_rec_nondata_replace_occured <= main_rtio_core_outputs_record17_rec_nondata_replace_occured;
			main_rtio_core_outputs_record29_rec_payload_channel <= main_rtio_core_outputs_record17_rec_payload_channel;
			main_rtio_core_outputs_record29_rec_payload_fine_ts <= main_rtio_core_outputs_record17_rec_payload_fine_ts;
			main_rtio_core_outputs_record29_rec_payload_address <= main_rtio_core_outputs_record17_rec_payload_address;
			main_rtio_core_outputs_record29_rec_payload_data <= main_rtio_core_outputs_record17_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record18_rec_valid), main_rtio_core_outputs_record18_rec_payload_channel} == {(~main_rtio_core_outputs_record22_rec_valid), main_rtio_core_outputs_record22_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record18_rec_seqn[10] == main_rtio_core_outputs_record18_rec_seqn[11]) & (main_rtio_core_outputs_record22_rec_seqn[10] == main_rtio_core_outputs_record22_rec_seqn[11])) & (main_rtio_core_outputs_record18_rec_seqn[11] != main_rtio_core_outputs_record22_rec_seqn[11])) ? main_rtio_core_outputs_record18_rec_seqn[11] : (main_rtio_core_outputs_record18_rec_seqn < main_rtio_core_outputs_record22_rec_seqn))) begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
		end
		main_rtio_core_outputs_record26_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference12;
		main_rtio_core_outputs_record30_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record18_rec_valid), main_rtio_core_outputs_record18_rec_payload_channel} < {(~main_rtio_core_outputs_record22_rec_valid), main_rtio_core_outputs_record22_rec_payload_channel})) begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record26_rec_valid <= main_rtio_core_outputs_record22_rec_valid;
			main_rtio_core_outputs_record26_rec_seqn <= main_rtio_core_outputs_record22_rec_seqn;
			main_rtio_core_outputs_record26_rec_replace_occured <= main_rtio_core_outputs_record22_rec_replace_occured;
			main_rtio_core_outputs_record26_rec_nondata_replace_occured <= main_rtio_core_outputs_record22_rec_nondata_replace_occured;
			main_rtio_core_outputs_record26_rec_payload_channel <= main_rtio_core_outputs_record22_rec_payload_channel;
			main_rtio_core_outputs_record26_rec_payload_fine_ts <= main_rtio_core_outputs_record22_rec_payload_fine_ts;
			main_rtio_core_outputs_record26_rec_payload_address <= main_rtio_core_outputs_record22_rec_payload_address;
			main_rtio_core_outputs_record26_rec_payload_data <= main_rtio_core_outputs_record22_rec_payload_data;
			main_rtio_core_outputs_record30_rec_valid <= main_rtio_core_outputs_record18_rec_valid;
			main_rtio_core_outputs_record30_rec_seqn <= main_rtio_core_outputs_record18_rec_seqn;
			main_rtio_core_outputs_record30_rec_replace_occured <= main_rtio_core_outputs_record18_rec_replace_occured;
			main_rtio_core_outputs_record30_rec_nondata_replace_occured <= main_rtio_core_outputs_record18_rec_nondata_replace_occured;
			main_rtio_core_outputs_record30_rec_payload_channel <= main_rtio_core_outputs_record18_rec_payload_channel;
			main_rtio_core_outputs_record30_rec_payload_fine_ts <= main_rtio_core_outputs_record18_rec_payload_fine_ts;
			main_rtio_core_outputs_record30_rec_payload_address <= main_rtio_core_outputs_record18_rec_payload_address;
			main_rtio_core_outputs_record30_rec_payload_data <= main_rtio_core_outputs_record18_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record19_rec_valid), main_rtio_core_outputs_record19_rec_payload_channel} == {(~main_rtio_core_outputs_record23_rec_valid), main_rtio_core_outputs_record23_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record19_rec_seqn[10] == main_rtio_core_outputs_record19_rec_seqn[11]) & (main_rtio_core_outputs_record23_rec_seqn[10] == main_rtio_core_outputs_record23_rec_seqn[11])) & (main_rtio_core_outputs_record19_rec_seqn[11] != main_rtio_core_outputs_record23_rec_seqn[11])) ? main_rtio_core_outputs_record19_rec_seqn[11] : (main_rtio_core_outputs_record19_rec_seqn < main_rtio_core_outputs_record23_rec_seqn))) begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
		end
		main_rtio_core_outputs_record27_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference13;
		main_rtio_core_outputs_record31_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record19_rec_valid), main_rtio_core_outputs_record19_rec_payload_channel} < {(~main_rtio_core_outputs_record23_rec_valid), main_rtio_core_outputs_record23_rec_payload_channel})) begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record27_rec_valid <= main_rtio_core_outputs_record23_rec_valid;
			main_rtio_core_outputs_record27_rec_seqn <= main_rtio_core_outputs_record23_rec_seqn;
			main_rtio_core_outputs_record27_rec_replace_occured <= main_rtio_core_outputs_record23_rec_replace_occured;
			main_rtio_core_outputs_record27_rec_nondata_replace_occured <= main_rtio_core_outputs_record23_rec_nondata_replace_occured;
			main_rtio_core_outputs_record27_rec_payload_channel <= main_rtio_core_outputs_record23_rec_payload_channel;
			main_rtio_core_outputs_record27_rec_payload_fine_ts <= main_rtio_core_outputs_record23_rec_payload_fine_ts;
			main_rtio_core_outputs_record27_rec_payload_address <= main_rtio_core_outputs_record23_rec_payload_address;
			main_rtio_core_outputs_record27_rec_payload_data <= main_rtio_core_outputs_record23_rec_payload_data;
			main_rtio_core_outputs_record31_rec_valid <= main_rtio_core_outputs_record19_rec_valid;
			main_rtio_core_outputs_record31_rec_seqn <= main_rtio_core_outputs_record19_rec_seqn;
			main_rtio_core_outputs_record31_rec_replace_occured <= main_rtio_core_outputs_record19_rec_replace_occured;
			main_rtio_core_outputs_record31_rec_nondata_replace_occured <= main_rtio_core_outputs_record19_rec_nondata_replace_occured;
			main_rtio_core_outputs_record31_rec_payload_channel <= main_rtio_core_outputs_record19_rec_payload_channel;
			main_rtio_core_outputs_record31_rec_payload_fine_ts <= main_rtio_core_outputs_record19_rec_payload_fine_ts;
			main_rtio_core_outputs_record31_rec_payload_address <= main_rtio_core_outputs_record19_rec_payload_address;
			main_rtio_core_outputs_record31_rec_payload_data <= main_rtio_core_outputs_record19_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record26_rec_valid), main_rtio_core_outputs_record26_rec_payload_channel} == {(~main_rtio_core_outputs_record28_rec_valid), main_rtio_core_outputs_record28_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record26_rec_seqn[10] == main_rtio_core_outputs_record26_rec_seqn[11]) & (main_rtio_core_outputs_record28_rec_seqn[10] == main_rtio_core_outputs_record28_rec_seqn[11])) & (main_rtio_core_outputs_record26_rec_seqn[11] != main_rtio_core_outputs_record28_rec_seqn[11])) ? main_rtio_core_outputs_record26_rec_seqn[11] : (main_rtio_core_outputs_record26_rec_seqn < main_rtio_core_outputs_record28_rec_seqn))) begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
		end
		main_rtio_core_outputs_record34_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference14;
		main_rtio_core_outputs_record36_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record26_rec_valid), main_rtio_core_outputs_record26_rec_payload_channel} < {(~main_rtio_core_outputs_record28_rec_valid), main_rtio_core_outputs_record28_rec_payload_channel})) begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record34_rec_valid <= main_rtio_core_outputs_record28_rec_valid;
			main_rtio_core_outputs_record34_rec_seqn <= main_rtio_core_outputs_record28_rec_seqn;
			main_rtio_core_outputs_record34_rec_replace_occured <= main_rtio_core_outputs_record28_rec_replace_occured;
			main_rtio_core_outputs_record34_rec_nondata_replace_occured <= main_rtio_core_outputs_record28_rec_nondata_replace_occured;
			main_rtio_core_outputs_record34_rec_payload_channel <= main_rtio_core_outputs_record28_rec_payload_channel;
			main_rtio_core_outputs_record34_rec_payload_fine_ts <= main_rtio_core_outputs_record28_rec_payload_fine_ts;
			main_rtio_core_outputs_record34_rec_payload_address <= main_rtio_core_outputs_record28_rec_payload_address;
			main_rtio_core_outputs_record34_rec_payload_data <= main_rtio_core_outputs_record28_rec_payload_data;
			main_rtio_core_outputs_record36_rec_valid <= main_rtio_core_outputs_record26_rec_valid;
			main_rtio_core_outputs_record36_rec_seqn <= main_rtio_core_outputs_record26_rec_seqn;
			main_rtio_core_outputs_record36_rec_replace_occured <= main_rtio_core_outputs_record26_rec_replace_occured;
			main_rtio_core_outputs_record36_rec_nondata_replace_occured <= main_rtio_core_outputs_record26_rec_nondata_replace_occured;
			main_rtio_core_outputs_record36_rec_payload_channel <= main_rtio_core_outputs_record26_rec_payload_channel;
			main_rtio_core_outputs_record36_rec_payload_fine_ts <= main_rtio_core_outputs_record26_rec_payload_fine_ts;
			main_rtio_core_outputs_record36_rec_payload_address <= main_rtio_core_outputs_record26_rec_payload_address;
			main_rtio_core_outputs_record36_rec_payload_data <= main_rtio_core_outputs_record26_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record27_rec_valid), main_rtio_core_outputs_record27_rec_payload_channel} == {(~main_rtio_core_outputs_record29_rec_valid), main_rtio_core_outputs_record29_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record27_rec_seqn[10] == main_rtio_core_outputs_record27_rec_seqn[11]) & (main_rtio_core_outputs_record29_rec_seqn[10] == main_rtio_core_outputs_record29_rec_seqn[11])) & (main_rtio_core_outputs_record27_rec_seqn[11] != main_rtio_core_outputs_record29_rec_seqn[11])) ? main_rtio_core_outputs_record27_rec_seqn[11] : (main_rtio_core_outputs_record27_rec_seqn < main_rtio_core_outputs_record29_rec_seqn))) begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
		end
		main_rtio_core_outputs_record35_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference15;
		main_rtio_core_outputs_record37_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record27_rec_valid), main_rtio_core_outputs_record27_rec_payload_channel} < {(~main_rtio_core_outputs_record29_rec_valid), main_rtio_core_outputs_record29_rec_payload_channel})) begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record35_rec_valid <= main_rtio_core_outputs_record29_rec_valid;
			main_rtio_core_outputs_record35_rec_seqn <= main_rtio_core_outputs_record29_rec_seqn;
			main_rtio_core_outputs_record35_rec_replace_occured <= main_rtio_core_outputs_record29_rec_replace_occured;
			main_rtio_core_outputs_record35_rec_nondata_replace_occured <= main_rtio_core_outputs_record29_rec_nondata_replace_occured;
			main_rtio_core_outputs_record35_rec_payload_channel <= main_rtio_core_outputs_record29_rec_payload_channel;
			main_rtio_core_outputs_record35_rec_payload_fine_ts <= main_rtio_core_outputs_record29_rec_payload_fine_ts;
			main_rtio_core_outputs_record35_rec_payload_address <= main_rtio_core_outputs_record29_rec_payload_address;
			main_rtio_core_outputs_record35_rec_payload_data <= main_rtio_core_outputs_record29_rec_payload_data;
			main_rtio_core_outputs_record37_rec_valid <= main_rtio_core_outputs_record27_rec_valid;
			main_rtio_core_outputs_record37_rec_seqn <= main_rtio_core_outputs_record27_rec_seqn;
			main_rtio_core_outputs_record37_rec_replace_occured <= main_rtio_core_outputs_record27_rec_replace_occured;
			main_rtio_core_outputs_record37_rec_nondata_replace_occured <= main_rtio_core_outputs_record27_rec_nondata_replace_occured;
			main_rtio_core_outputs_record37_rec_payload_channel <= main_rtio_core_outputs_record27_rec_payload_channel;
			main_rtio_core_outputs_record37_rec_payload_fine_ts <= main_rtio_core_outputs_record27_rec_payload_fine_ts;
			main_rtio_core_outputs_record37_rec_payload_address <= main_rtio_core_outputs_record27_rec_payload_address;
			main_rtio_core_outputs_record37_rec_payload_data <= main_rtio_core_outputs_record27_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record32_rec_valid <= main_rtio_core_outputs_record24_rec_valid;
	main_rtio_core_outputs_record32_rec_seqn <= main_rtio_core_outputs_record24_rec_seqn;
	main_rtio_core_outputs_record32_rec_replace_occured <= main_rtio_core_outputs_record24_rec_replace_occured;
	main_rtio_core_outputs_record32_rec_nondata_replace_occured <= main_rtio_core_outputs_record24_rec_nondata_replace_occured;
	main_rtio_core_outputs_record32_rec_payload_channel <= main_rtio_core_outputs_record24_rec_payload_channel;
	main_rtio_core_outputs_record32_rec_payload_fine_ts <= main_rtio_core_outputs_record24_rec_payload_fine_ts;
	main_rtio_core_outputs_record32_rec_payload_address <= main_rtio_core_outputs_record24_rec_payload_address;
	main_rtio_core_outputs_record32_rec_payload_data <= main_rtio_core_outputs_record24_rec_payload_data;
	main_rtio_core_outputs_record33_rec_valid <= main_rtio_core_outputs_record25_rec_valid;
	main_rtio_core_outputs_record33_rec_seqn <= main_rtio_core_outputs_record25_rec_seqn;
	main_rtio_core_outputs_record33_rec_replace_occured <= main_rtio_core_outputs_record25_rec_replace_occured;
	main_rtio_core_outputs_record33_rec_nondata_replace_occured <= main_rtio_core_outputs_record25_rec_nondata_replace_occured;
	main_rtio_core_outputs_record33_rec_payload_channel <= main_rtio_core_outputs_record25_rec_payload_channel;
	main_rtio_core_outputs_record33_rec_payload_fine_ts <= main_rtio_core_outputs_record25_rec_payload_fine_ts;
	main_rtio_core_outputs_record33_rec_payload_address <= main_rtio_core_outputs_record25_rec_payload_address;
	main_rtio_core_outputs_record33_rec_payload_data <= main_rtio_core_outputs_record25_rec_payload_data;
	main_rtio_core_outputs_record38_rec_valid <= main_rtio_core_outputs_record30_rec_valid;
	main_rtio_core_outputs_record38_rec_seqn <= main_rtio_core_outputs_record30_rec_seqn;
	main_rtio_core_outputs_record38_rec_replace_occured <= main_rtio_core_outputs_record30_rec_replace_occured;
	main_rtio_core_outputs_record38_rec_nondata_replace_occured <= main_rtio_core_outputs_record30_rec_nondata_replace_occured;
	main_rtio_core_outputs_record38_rec_payload_channel <= main_rtio_core_outputs_record30_rec_payload_channel;
	main_rtio_core_outputs_record38_rec_payload_fine_ts <= main_rtio_core_outputs_record30_rec_payload_fine_ts;
	main_rtio_core_outputs_record38_rec_payload_address <= main_rtio_core_outputs_record30_rec_payload_address;
	main_rtio_core_outputs_record38_rec_payload_data <= main_rtio_core_outputs_record30_rec_payload_data;
	main_rtio_core_outputs_record39_rec_valid <= main_rtio_core_outputs_record31_rec_valid;
	main_rtio_core_outputs_record39_rec_seqn <= main_rtio_core_outputs_record31_rec_seqn;
	main_rtio_core_outputs_record39_rec_replace_occured <= main_rtio_core_outputs_record31_rec_replace_occured;
	main_rtio_core_outputs_record39_rec_nondata_replace_occured <= main_rtio_core_outputs_record31_rec_nondata_replace_occured;
	main_rtio_core_outputs_record39_rec_payload_channel <= main_rtio_core_outputs_record31_rec_payload_channel;
	main_rtio_core_outputs_record39_rec_payload_fine_ts <= main_rtio_core_outputs_record31_rec_payload_fine_ts;
	main_rtio_core_outputs_record39_rec_payload_address <= main_rtio_core_outputs_record31_rec_payload_address;
	main_rtio_core_outputs_record39_rec_payload_data <= main_rtio_core_outputs_record31_rec_payload_data;
	if (({(~main_rtio_core_outputs_record33_rec_valid), main_rtio_core_outputs_record33_rec_payload_channel} == {(~main_rtio_core_outputs_record34_rec_valid), main_rtio_core_outputs_record34_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record33_rec_seqn[10] == main_rtio_core_outputs_record33_rec_seqn[11]) & (main_rtio_core_outputs_record34_rec_seqn[10] == main_rtio_core_outputs_record34_rec_seqn[11])) & (main_rtio_core_outputs_record33_rec_seqn[11] != main_rtio_core_outputs_record34_rec_seqn[11])) ? main_rtio_core_outputs_record33_rec_seqn[11] : (main_rtio_core_outputs_record33_rec_seqn < main_rtio_core_outputs_record34_rec_seqn))) begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
		end
		main_rtio_core_outputs_record41_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference16;
		main_rtio_core_outputs_record42_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record33_rec_valid), main_rtio_core_outputs_record33_rec_payload_channel} < {(~main_rtio_core_outputs_record34_rec_valid), main_rtio_core_outputs_record34_rec_payload_channel})) begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record41_rec_valid <= main_rtio_core_outputs_record34_rec_valid;
			main_rtio_core_outputs_record41_rec_seqn <= main_rtio_core_outputs_record34_rec_seqn;
			main_rtio_core_outputs_record41_rec_replace_occured <= main_rtio_core_outputs_record34_rec_replace_occured;
			main_rtio_core_outputs_record41_rec_nondata_replace_occured <= main_rtio_core_outputs_record34_rec_nondata_replace_occured;
			main_rtio_core_outputs_record41_rec_payload_channel <= main_rtio_core_outputs_record34_rec_payload_channel;
			main_rtio_core_outputs_record41_rec_payload_fine_ts <= main_rtio_core_outputs_record34_rec_payload_fine_ts;
			main_rtio_core_outputs_record41_rec_payload_address <= main_rtio_core_outputs_record34_rec_payload_address;
			main_rtio_core_outputs_record41_rec_payload_data <= main_rtio_core_outputs_record34_rec_payload_data;
			main_rtio_core_outputs_record42_rec_valid <= main_rtio_core_outputs_record33_rec_valid;
			main_rtio_core_outputs_record42_rec_seqn <= main_rtio_core_outputs_record33_rec_seqn;
			main_rtio_core_outputs_record42_rec_replace_occured <= main_rtio_core_outputs_record33_rec_replace_occured;
			main_rtio_core_outputs_record42_rec_nondata_replace_occured <= main_rtio_core_outputs_record33_rec_nondata_replace_occured;
			main_rtio_core_outputs_record42_rec_payload_channel <= main_rtio_core_outputs_record33_rec_payload_channel;
			main_rtio_core_outputs_record42_rec_payload_fine_ts <= main_rtio_core_outputs_record33_rec_payload_fine_ts;
			main_rtio_core_outputs_record42_rec_payload_address <= main_rtio_core_outputs_record33_rec_payload_address;
			main_rtio_core_outputs_record42_rec_payload_data <= main_rtio_core_outputs_record33_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record35_rec_valid), main_rtio_core_outputs_record35_rec_payload_channel} == {(~main_rtio_core_outputs_record36_rec_valid), main_rtio_core_outputs_record36_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record35_rec_seqn[10] == main_rtio_core_outputs_record35_rec_seqn[11]) & (main_rtio_core_outputs_record36_rec_seqn[10] == main_rtio_core_outputs_record36_rec_seqn[11])) & (main_rtio_core_outputs_record35_rec_seqn[11] != main_rtio_core_outputs_record36_rec_seqn[11])) ? main_rtio_core_outputs_record35_rec_seqn[11] : (main_rtio_core_outputs_record35_rec_seqn < main_rtio_core_outputs_record36_rec_seqn))) begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
		end
		main_rtio_core_outputs_record43_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference17;
		main_rtio_core_outputs_record44_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record35_rec_valid), main_rtio_core_outputs_record35_rec_payload_channel} < {(~main_rtio_core_outputs_record36_rec_valid), main_rtio_core_outputs_record36_rec_payload_channel})) begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record43_rec_valid <= main_rtio_core_outputs_record36_rec_valid;
			main_rtio_core_outputs_record43_rec_seqn <= main_rtio_core_outputs_record36_rec_seqn;
			main_rtio_core_outputs_record43_rec_replace_occured <= main_rtio_core_outputs_record36_rec_replace_occured;
			main_rtio_core_outputs_record43_rec_nondata_replace_occured <= main_rtio_core_outputs_record36_rec_nondata_replace_occured;
			main_rtio_core_outputs_record43_rec_payload_channel <= main_rtio_core_outputs_record36_rec_payload_channel;
			main_rtio_core_outputs_record43_rec_payload_fine_ts <= main_rtio_core_outputs_record36_rec_payload_fine_ts;
			main_rtio_core_outputs_record43_rec_payload_address <= main_rtio_core_outputs_record36_rec_payload_address;
			main_rtio_core_outputs_record43_rec_payload_data <= main_rtio_core_outputs_record36_rec_payload_data;
			main_rtio_core_outputs_record44_rec_valid <= main_rtio_core_outputs_record35_rec_valid;
			main_rtio_core_outputs_record44_rec_seqn <= main_rtio_core_outputs_record35_rec_seqn;
			main_rtio_core_outputs_record44_rec_replace_occured <= main_rtio_core_outputs_record35_rec_replace_occured;
			main_rtio_core_outputs_record44_rec_nondata_replace_occured <= main_rtio_core_outputs_record35_rec_nondata_replace_occured;
			main_rtio_core_outputs_record44_rec_payload_channel <= main_rtio_core_outputs_record35_rec_payload_channel;
			main_rtio_core_outputs_record44_rec_payload_fine_ts <= main_rtio_core_outputs_record35_rec_payload_fine_ts;
			main_rtio_core_outputs_record44_rec_payload_address <= main_rtio_core_outputs_record35_rec_payload_address;
			main_rtio_core_outputs_record44_rec_payload_data <= main_rtio_core_outputs_record35_rec_payload_data;
		end
	end
	if (({(~main_rtio_core_outputs_record37_rec_valid), main_rtio_core_outputs_record37_rec_payload_channel} == {(~main_rtio_core_outputs_record38_rec_valid), main_rtio_core_outputs_record38_rec_payload_channel})) begin
		if (((((main_rtio_core_outputs_record37_rec_seqn[10] == main_rtio_core_outputs_record37_rec_seqn[11]) & (main_rtio_core_outputs_record38_rec_seqn[10] == main_rtio_core_outputs_record38_rec_seqn[11])) & (main_rtio_core_outputs_record37_rec_seqn[11] != main_rtio_core_outputs_record38_rec_seqn[11])) ? main_rtio_core_outputs_record37_rec_seqn[11] : (main_rtio_core_outputs_record37_rec_seqn < main_rtio_core_outputs_record38_rec_seqn))) begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
		end
		main_rtio_core_outputs_record45_rec_replace_occured <= 1'd1;
		main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_nondata_difference18;
		main_rtio_core_outputs_record46_rec_valid <= 1'd0;
	end else begin
		if (({(~main_rtio_core_outputs_record37_rec_valid), main_rtio_core_outputs_record37_rec_payload_channel} < {(~main_rtio_core_outputs_record38_rec_valid), main_rtio_core_outputs_record38_rec_payload_channel})) begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
		end else begin
			main_rtio_core_outputs_record45_rec_valid <= main_rtio_core_outputs_record38_rec_valid;
			main_rtio_core_outputs_record45_rec_seqn <= main_rtio_core_outputs_record38_rec_seqn;
			main_rtio_core_outputs_record45_rec_replace_occured <= main_rtio_core_outputs_record38_rec_replace_occured;
			main_rtio_core_outputs_record45_rec_nondata_replace_occured <= main_rtio_core_outputs_record38_rec_nondata_replace_occured;
			main_rtio_core_outputs_record45_rec_payload_channel <= main_rtio_core_outputs_record38_rec_payload_channel;
			main_rtio_core_outputs_record45_rec_payload_fine_ts <= main_rtio_core_outputs_record38_rec_payload_fine_ts;
			main_rtio_core_outputs_record45_rec_payload_address <= main_rtio_core_outputs_record38_rec_payload_address;
			main_rtio_core_outputs_record45_rec_payload_data <= main_rtio_core_outputs_record38_rec_payload_data;
			main_rtio_core_outputs_record46_rec_valid <= main_rtio_core_outputs_record37_rec_valid;
			main_rtio_core_outputs_record46_rec_seqn <= main_rtio_core_outputs_record37_rec_seqn;
			main_rtio_core_outputs_record46_rec_replace_occured <= main_rtio_core_outputs_record37_rec_replace_occured;
			main_rtio_core_outputs_record46_rec_nondata_replace_occured <= main_rtio_core_outputs_record37_rec_nondata_replace_occured;
			main_rtio_core_outputs_record46_rec_payload_channel <= main_rtio_core_outputs_record37_rec_payload_channel;
			main_rtio_core_outputs_record46_rec_payload_fine_ts <= main_rtio_core_outputs_record37_rec_payload_fine_ts;
			main_rtio_core_outputs_record46_rec_payload_address <= main_rtio_core_outputs_record37_rec_payload_address;
			main_rtio_core_outputs_record46_rec_payload_data <= main_rtio_core_outputs_record37_rec_payload_data;
		end
	end
	main_rtio_core_outputs_record40_rec_valid <= main_rtio_core_outputs_record32_rec_valid;
	main_rtio_core_outputs_record40_rec_seqn <= main_rtio_core_outputs_record32_rec_seqn;
	main_rtio_core_outputs_record40_rec_replace_occured <= main_rtio_core_outputs_record32_rec_replace_occured;
	main_rtio_core_outputs_record40_rec_nondata_replace_occured <= main_rtio_core_outputs_record32_rec_nondata_replace_occured;
	main_rtio_core_outputs_record40_rec_payload_channel <= main_rtio_core_outputs_record32_rec_payload_channel;
	main_rtio_core_outputs_record40_rec_payload_fine_ts <= main_rtio_core_outputs_record32_rec_payload_fine_ts;
	main_rtio_core_outputs_record40_rec_payload_address <= main_rtio_core_outputs_record32_rec_payload_address;
	main_rtio_core_outputs_record40_rec_payload_data <= main_rtio_core_outputs_record32_rec_payload_data;
	main_rtio_core_outputs_record47_rec_valid <= main_rtio_core_outputs_record39_rec_valid;
	main_rtio_core_outputs_record47_rec_seqn <= main_rtio_core_outputs_record39_rec_seqn;
	main_rtio_core_outputs_record47_rec_replace_occured <= main_rtio_core_outputs_record39_rec_replace_occured;
	main_rtio_core_outputs_record47_rec_nondata_replace_occured <= main_rtio_core_outputs_record39_rec_nondata_replace_occured;
	main_rtio_core_outputs_record47_rec_payload_channel <= main_rtio_core_outputs_record39_rec_payload_channel;
	main_rtio_core_outputs_record47_rec_payload_fine_ts <= main_rtio_core_outputs_record39_rec_payload_fine_ts;
	main_rtio_core_outputs_record47_rec_payload_address <= main_rtio_core_outputs_record39_rec_payload_address;
	main_rtio_core_outputs_record47_rec_payload_data <= main_rtio_core_outputs_record39_rec_payload_data;
	main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_next_binary;
	main_rtio_core_inputs_asyncfifo0_graycounter0_q <= main_rtio_core_inputs_asyncfifo0_graycounter0_q_next;
	if (main_rtio_core_inputs_blindtransfer0_i) begin
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer0_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer0_ps_i) begin
		main_rtio_core_inputs_blindtransfer0_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer0_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_next_binary;
	main_rtio_core_inputs_asyncfifo1_graycounter2_q <= main_rtio_core_inputs_asyncfifo1_graycounter2_q_next;
	if (main_rtio_core_inputs_blindtransfer1_i) begin
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer1_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer1_ps_i) begin
		main_rtio_core_inputs_blindtransfer1_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer1_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_next_binary;
	main_rtio_core_inputs_asyncfifo2_graycounter4_q <= main_rtio_core_inputs_asyncfifo2_graycounter4_q_next;
	if (main_rtio_core_inputs_blindtransfer2_i) begin
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer2_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer2_ps_i) begin
		main_rtio_core_inputs_blindtransfer2_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer2_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_next_binary;
	main_rtio_core_inputs_asyncfifo3_graycounter6_q <= main_rtio_core_inputs_asyncfifo3_graycounter6_q_next;
	if (main_rtio_core_inputs_blindtransfer3_i) begin
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer3_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer3_ps_i) begin
		main_rtio_core_inputs_blindtransfer3_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer3_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_next_binary;
	main_rtio_core_inputs_asyncfifo4_graycounter8_q <= main_rtio_core_inputs_asyncfifo4_graycounter8_q_next;
	if (main_rtio_core_inputs_blindtransfer4_i) begin
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer4_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer4_ps_i) begin
		main_rtio_core_inputs_blindtransfer4_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer4_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_next_binary;
	main_rtio_core_inputs_asyncfifo5_graycounter10_q <= main_rtio_core_inputs_asyncfifo5_graycounter10_q_next;
	if (main_rtio_core_inputs_blindtransfer5_i) begin
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer5_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer5_ps_i) begin
		main_rtio_core_inputs_blindtransfer5_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer5_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_next_binary;
	main_rtio_core_inputs_asyncfifo6_graycounter12_q <= main_rtio_core_inputs_asyncfifo6_graycounter12_q_next;
	if (main_rtio_core_inputs_blindtransfer6_i) begin
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer6_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer6_ps_i) begin
		main_rtio_core_inputs_blindtransfer6_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer6_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_next_binary;
	main_rtio_core_inputs_asyncfifo7_graycounter14_q <= main_rtio_core_inputs_asyncfifo7_graycounter14_q_next;
	if (main_rtio_core_inputs_blindtransfer7_i) begin
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer7_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer7_ps_i) begin
		main_rtio_core_inputs_blindtransfer7_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer7_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_next_binary;
	main_rtio_core_inputs_asyncfifo8_graycounter16_q <= main_rtio_core_inputs_asyncfifo8_graycounter16_q_next;
	if (main_rtio_core_inputs_blindtransfer8_i) begin
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer8_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer8_ps_i) begin
		main_rtio_core_inputs_blindtransfer8_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer8_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_next_binary;
	main_rtio_core_inputs_asyncfifo9_graycounter18_q <= main_rtio_core_inputs_asyncfifo9_graycounter18_q_next;
	if (main_rtio_core_inputs_blindtransfer9_i) begin
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer9_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer9_ps_i) begin
		main_rtio_core_inputs_blindtransfer9_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer9_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_next_binary;
	main_rtio_core_inputs_asyncfifo10_graycounter20_q <= main_rtio_core_inputs_asyncfifo10_graycounter20_q_next;
	if (main_rtio_core_inputs_blindtransfer10_i) begin
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer10_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer10_ps_i) begin
		main_rtio_core_inputs_blindtransfer10_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer10_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_o;
	main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary <= main_rtio_core_inputs_asyncfifo11_graycounter22_q_next_binary;
	main_rtio_core_inputs_asyncfifo11_graycounter22_q <= main_rtio_core_inputs_asyncfifo11_graycounter22_q_next;
	if (main_rtio_core_inputs_blindtransfer11_i) begin
		main_rtio_core_inputs_blindtransfer11_blind <= 1'd1;
	end
	if (main_rtio_core_inputs_blindtransfer11_ps_ack_o) begin
		main_rtio_core_inputs_blindtransfer11_blind <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer11_ps_i) begin
		main_rtio_core_inputs_blindtransfer11_ps_toggle_i <= (~main_rtio_core_inputs_blindtransfer11_ps_toggle_i);
	end
	main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o_r <= main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_o;
	if (main_rtio_core_o_collision_sync_i) begin
		main_rtio_core_o_collision_sync_blind <= 1'd1;
	end
	if (main_rtio_core_o_collision_sync_ps_ack_o) begin
		main_rtio_core_o_collision_sync_blind <= 1'd0;
	end
	if (main_rtio_core_o_collision_sync_ps_i) begin
		main_rtio_core_o_collision_sync_bxfer_data <= main_rtio_core_o_collision_sync_data_i;
	end
	if (main_rtio_core_o_collision_sync_ps_i) begin
		main_rtio_core_o_collision_sync_ps_toggle_i <= (~main_rtio_core_o_collision_sync_ps_toggle_i);
	end
	main_rtio_core_o_collision_sync_ps_ack_toggle_o_r <= main_rtio_core_o_collision_sync_ps_ack_toggle_o;
	if (main_rtio_core_o_busy_sync_i) begin
		main_rtio_core_o_busy_sync_blind <= 1'd1;
	end
	if (main_rtio_core_o_busy_sync_ps_ack_o) begin
		main_rtio_core_o_busy_sync_blind <= 1'd0;
	end
	if (main_rtio_core_o_busy_sync_ps_i) begin
		main_rtio_core_o_busy_sync_bxfer_data <= main_rtio_core_o_busy_sync_data_i;
	end
	if (main_rtio_core_o_busy_sync_ps_i) begin
		main_rtio_core_o_busy_sync_ps_toggle_i <= (~main_rtio_core_o_busy_sync_ps_toggle_i);
	end
	main_rtio_core_o_busy_sync_ps_ack_toggle_o_r <= main_rtio_core_o_busy_sync_ps_ack_toggle_o;
	main_mon_bussynchronizer28_starter <= 1'd0;
	if (main_mon_bussynchronizer28_pong_o) begin
		main_mon_bussynchronizer28_ibuffer <= main_mon_bussynchronizer28_i;
	end
	if (main_mon_bussynchronizer28_ping_i) begin
		main_mon_bussynchronizer28_ping_toggle_i <= (~main_mon_bussynchronizer28_ping_toggle_i);
	end
	main_mon_bussynchronizer28_pong_toggle_o_r <= main_mon_bussynchronizer28_pong_toggle_o;
	if (main_mon_bussynchronizer28_wait) begin
		if ((~main_mon_bussynchronizer28_done)) begin
			main_mon_bussynchronizer28_count <= (main_mon_bussynchronizer28_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer28_count <= 8'd128;
	end
	main_mon_bussynchronizer29_starter <= 1'd0;
	if (main_mon_bussynchronizer29_pong_o) begin
		main_mon_bussynchronizer29_ibuffer <= main_mon_bussynchronizer29_i;
	end
	if (main_mon_bussynchronizer29_ping_i) begin
		main_mon_bussynchronizer29_ping_toggle_i <= (~main_mon_bussynchronizer29_ping_toggle_i);
	end
	main_mon_bussynchronizer29_pong_toggle_o_r <= main_mon_bussynchronizer29_pong_toggle_o;
	if (main_mon_bussynchronizer29_wait) begin
		if ((~main_mon_bussynchronizer29_done)) begin
			main_mon_bussynchronizer29_count <= (main_mon_bussynchronizer29_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer29_count <= 8'd128;
	end
	main_mon_bussynchronizer30_starter <= 1'd0;
	if (main_mon_bussynchronizer30_pong_o) begin
		main_mon_bussynchronizer30_ibuffer <= main_mon_bussynchronizer30_i;
	end
	if (main_mon_bussynchronizer30_ping_i) begin
		main_mon_bussynchronizer30_ping_toggle_i <= (~main_mon_bussynchronizer30_ping_toggle_i);
	end
	main_mon_bussynchronizer30_pong_toggle_o_r <= main_mon_bussynchronizer30_pong_toggle_o;
	if (main_mon_bussynchronizer30_wait) begin
		if ((~main_mon_bussynchronizer30_done)) begin
			main_mon_bussynchronizer30_count <= (main_mon_bussynchronizer30_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer30_count <= 8'd128;
	end
	main_mon_bussynchronizer31_starter <= 1'd0;
	if (main_mon_bussynchronizer31_pong_o) begin
		main_mon_bussynchronizer31_ibuffer <= main_mon_bussynchronizer31_i;
	end
	if (main_mon_bussynchronizer31_ping_i) begin
		main_mon_bussynchronizer31_ping_toggle_i <= (~main_mon_bussynchronizer31_ping_toggle_i);
	end
	main_mon_bussynchronizer31_pong_toggle_o_r <= main_mon_bussynchronizer31_pong_toggle_o;
	if (main_mon_bussynchronizer31_wait) begin
		if ((~main_mon_bussynchronizer31_done)) begin
			main_mon_bussynchronizer31_count <= (main_mon_bussynchronizer31_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer31_count <= 8'd128;
	end
	main_mon_bussynchronizer32_starter <= 1'd0;
	if (main_mon_bussynchronizer32_pong_o) begin
		main_mon_bussynchronizer32_ibuffer <= main_mon_bussynchronizer32_i;
	end
	if (main_mon_bussynchronizer32_ping_i) begin
		main_mon_bussynchronizer32_ping_toggle_i <= (~main_mon_bussynchronizer32_ping_toggle_i);
	end
	main_mon_bussynchronizer32_pong_toggle_o_r <= main_mon_bussynchronizer32_pong_toggle_o;
	if (main_mon_bussynchronizer32_wait) begin
		if ((~main_mon_bussynchronizer32_done)) begin
			main_mon_bussynchronizer32_count <= (main_mon_bussynchronizer32_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer32_count <= 8'd128;
	end
	main_mon_bussynchronizer33_starter <= 1'd0;
	if (main_mon_bussynchronizer33_pong_o) begin
		main_mon_bussynchronizer33_ibuffer <= main_mon_bussynchronizer33_i;
	end
	if (main_mon_bussynchronizer33_ping_i) begin
		main_mon_bussynchronizer33_ping_toggle_i <= (~main_mon_bussynchronizer33_ping_toggle_i);
	end
	main_mon_bussynchronizer33_pong_toggle_o_r <= main_mon_bussynchronizer33_pong_toggle_o;
	if (main_mon_bussynchronizer33_wait) begin
		if ((~main_mon_bussynchronizer33_done)) begin
			main_mon_bussynchronizer33_count <= (main_mon_bussynchronizer33_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer33_count <= 8'd128;
	end
	main_mon_bussynchronizer34_starter <= 1'd0;
	if (main_mon_bussynchronizer34_pong_o) begin
		main_mon_bussynchronizer34_ibuffer <= main_mon_bussynchronizer34_i;
	end
	if (main_mon_bussynchronizer34_ping_i) begin
		main_mon_bussynchronizer34_ping_toggle_i <= (~main_mon_bussynchronizer34_ping_toggle_i);
	end
	main_mon_bussynchronizer34_pong_toggle_o_r <= main_mon_bussynchronizer34_pong_toggle_o;
	if (main_mon_bussynchronizer34_wait) begin
		if ((~main_mon_bussynchronizer34_done)) begin
			main_mon_bussynchronizer34_count <= (main_mon_bussynchronizer34_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer34_count <= 8'd128;
	end
	main_mon_bussynchronizer35_starter <= 1'd0;
	if (main_mon_bussynchronizer35_pong_o) begin
		main_mon_bussynchronizer35_ibuffer <= main_mon_bussynchronizer35_i;
	end
	if (main_mon_bussynchronizer35_ping_i) begin
		main_mon_bussynchronizer35_ping_toggle_i <= (~main_mon_bussynchronizer35_ping_toggle_i);
	end
	main_mon_bussynchronizer35_pong_toggle_o_r <= main_mon_bussynchronizer35_pong_toggle_o;
	if (main_mon_bussynchronizer35_wait) begin
		if ((~main_mon_bussynchronizer35_done)) begin
			main_mon_bussynchronizer35_count <= (main_mon_bussynchronizer35_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer35_count <= 8'd128;
	end
	main_mon_bussynchronizer36_starter <= 1'd0;
	if (main_mon_bussynchronizer36_pong_o) begin
		main_mon_bussynchronizer36_ibuffer <= main_mon_bussynchronizer36_i;
	end
	if (main_mon_bussynchronizer36_ping_i) begin
		main_mon_bussynchronizer36_ping_toggle_i <= (~main_mon_bussynchronizer36_ping_toggle_i);
	end
	main_mon_bussynchronizer36_pong_toggle_o_r <= main_mon_bussynchronizer36_pong_toggle_o;
	if (main_mon_bussynchronizer36_wait) begin
		if ((~main_mon_bussynchronizer36_done)) begin
			main_mon_bussynchronizer36_count <= (main_mon_bussynchronizer36_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer36_count <= 8'd128;
	end
	main_mon_bussynchronizer37_starter <= 1'd0;
	if (main_mon_bussynchronizer37_pong_o) begin
		main_mon_bussynchronizer37_ibuffer <= main_mon_bussynchronizer37_i;
	end
	if (main_mon_bussynchronizer37_ping_i) begin
		main_mon_bussynchronizer37_ping_toggle_i <= (~main_mon_bussynchronizer37_ping_toggle_i);
	end
	main_mon_bussynchronizer37_pong_toggle_o_r <= main_mon_bussynchronizer37_pong_toggle_o;
	if (main_mon_bussynchronizer37_wait) begin
		if ((~main_mon_bussynchronizer37_done)) begin
			main_mon_bussynchronizer37_count <= (main_mon_bussynchronizer37_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer37_count <= 8'd128;
	end
	main_mon_bussynchronizer38_starter <= 1'd0;
	if (main_mon_bussynchronizer38_pong_o) begin
		main_mon_bussynchronizer38_ibuffer <= main_mon_bussynchronizer38_i;
	end
	if (main_mon_bussynchronizer38_ping_i) begin
		main_mon_bussynchronizer38_ping_toggle_i <= (~main_mon_bussynchronizer38_ping_toggle_i);
	end
	main_mon_bussynchronizer38_pong_toggle_o_r <= main_mon_bussynchronizer38_pong_toggle_o;
	if (main_mon_bussynchronizer38_wait) begin
		if ((~main_mon_bussynchronizer38_done)) begin
			main_mon_bussynchronizer38_count <= (main_mon_bussynchronizer38_count - 1'd1);
		end
	end else begin
		main_mon_bussynchronizer38_count <= 8'd128;
	end
	if (rio_rst) begin
		main_output_8x0_stb <= 1'd0;
		main_output_8x1_stb <= 1'd0;
		main_output_8x2_stb <= 1'd0;
		main_inout_8x0_inout_8x0_ointerface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_sensitivity <= 2'd0;
		main_inout_8x0_inout_8x0_sample <= 1'd0;
		main_output_8x3_stb <= 1'd0;
		main_output_8x4_stb <= 1'd0;
		main_output_8x5_stb <= 1'd0;
		main_inout_8x1_inout_8x1_ointerface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_sensitivity <= 2'd0;
		main_inout_8x1_inout_8x1_sample <= 1'd0;
		main_output_8x6_stb <= 1'd0;
		main_output_8x7_stb <= 1'd0;
		main_output_8x8_stb <= 1'd0;
		main_inout_8x2_inout_8x2_ointerface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_sensitivity <= 2'd0;
		main_inout_8x2_inout_8x2_sample <= 1'd0;
		main_output_8x9_stb <= 1'd0;
		main_output_8x10_stb <= 1'd0;
		main_output_8x11_stb <= 1'd0;
		main_inout_8x3_inout_8x3_ointerface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_sensitivity <= 2'd0;
		main_inout_8x3_inout_8x3_sample <= 1'd0;
		main_inout_8x4_inout_8x4_ointerface4_stb <= 1'd0;
		main_inout_8x4_inout_8x4_sensitivity <= 2'd0;
		main_inout_8x4_inout_8x4_sample <= 1'd0;
		main_inout_8x5_inout_8x5_ointerface5_stb <= 1'd0;
		main_inout_8x5_inout_8x5_sensitivity <= 2'd0;
		main_inout_8x5_inout_8x5_sample <= 1'd0;
		main_inout_8x6_inout_8x6_ointerface6_stb <= 1'd0;
		main_inout_8x6_inout_8x6_sensitivity <= 2'd0;
		main_inout_8x6_inout_8x6_sample <= 1'd0;
		main_output0_stb <= 1'd0;
		main_output1_stb <= 1'd0;
		main_clockgen_stb <= 1'd0;
		main_clockgen_ftw <= 24'd0;
		main_spimaster0_ointerface0_stb <= 1'd0;
		main_spimaster1_ointerface1_stb <= 1'd0;
		main_spimaster2_ointerface2_stb <= 1'd0;
		main_spimaster3_ointerface3_stb <= 1'd0;
		main_spimaster4_ointerface4_stb <= 1'd0;
		main_ad9914_bus_adr <= 30'd0;
		main_ad9914_bus_dat_w <= 16'd0;
		main_ad9914_bus_sel <= 2'd0;
		main_ad9914_bus_we <= 1'd0;
		main_ad9914_stb <= 1'd0;
		main_ad9914_active <= 1'd0;
		main_ad9914_current_sel <= 15'd0;
		main_stb <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered0_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_readable <= 1'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q_binary <= 8'd0;
		main_rtio_core_outputs_gates_record0_valid <= 1'd0;
		main_rtio_core_outputs_gates_record1_valid <= 1'd0;
		main_rtio_core_outputs_gates_record2_valid <= 1'd0;
		main_rtio_core_outputs_gates_record3_valid <= 1'd0;
		main_rtio_core_outputs_gates_record4_valid <= 1'd0;
		main_rtio_core_outputs_gates_record5_valid <= 1'd0;
		main_rtio_core_outputs_gates_record6_valid <= 1'd0;
		main_rtio_core_outputs_gates_record7_valid <= 1'd0;
		main_rtio_core_outputs_collision <= 1'd0;
		main_rtio_core_outputs_busy <= 1'd0;
		main_rtio_core_outputs_record0_rec_valid <= 1'd0;
		main_rtio_core_outputs_record1_rec_valid <= 1'd0;
		main_rtio_core_outputs_record2_rec_valid <= 1'd0;
		main_rtio_core_outputs_record3_rec_valid <= 1'd0;
		main_rtio_core_outputs_record4_rec_valid <= 1'd0;
		main_rtio_core_outputs_record5_rec_valid <= 1'd0;
		main_rtio_core_outputs_record6_rec_valid <= 1'd0;
		main_rtio_core_outputs_record7_rec_valid <= 1'd0;
		main_rtio_core_outputs_record8_rec_valid <= 1'd0;
		main_rtio_core_outputs_record9_rec_valid <= 1'd0;
		main_rtio_core_outputs_record10_rec_valid <= 1'd0;
		main_rtio_core_outputs_record11_rec_valid <= 1'd0;
		main_rtio_core_outputs_record12_rec_valid <= 1'd0;
		main_rtio_core_outputs_record13_rec_valid <= 1'd0;
		main_rtio_core_outputs_record14_rec_valid <= 1'd0;
		main_rtio_core_outputs_record15_rec_valid <= 1'd0;
		main_rtio_core_outputs_record16_rec_valid <= 1'd0;
		main_rtio_core_outputs_record17_rec_valid <= 1'd0;
		main_rtio_core_outputs_record18_rec_valid <= 1'd0;
		main_rtio_core_outputs_record19_rec_valid <= 1'd0;
		main_rtio_core_outputs_record20_rec_valid <= 1'd0;
		main_rtio_core_outputs_record21_rec_valid <= 1'd0;
		main_rtio_core_outputs_record22_rec_valid <= 1'd0;
		main_rtio_core_outputs_record23_rec_valid <= 1'd0;
		main_rtio_core_outputs_record24_rec_valid <= 1'd0;
		main_rtio_core_outputs_record25_rec_valid <= 1'd0;
		main_rtio_core_outputs_record26_rec_valid <= 1'd0;
		main_rtio_core_outputs_record27_rec_valid <= 1'd0;
		main_rtio_core_outputs_record28_rec_valid <= 1'd0;
		main_rtio_core_outputs_record29_rec_valid <= 1'd0;
		main_rtio_core_outputs_record30_rec_valid <= 1'd0;
		main_rtio_core_outputs_record31_rec_valid <= 1'd0;
		main_rtio_core_outputs_record32_rec_valid <= 1'd0;
		main_rtio_core_outputs_record33_rec_valid <= 1'd0;
		main_rtio_core_outputs_record34_rec_valid <= 1'd0;
		main_rtio_core_outputs_record35_rec_valid <= 1'd0;
		main_rtio_core_outputs_record36_rec_valid <= 1'd0;
		main_rtio_core_outputs_record37_rec_valid <= 1'd0;
		main_rtio_core_outputs_record38_rec_valid <= 1'd0;
		main_rtio_core_outputs_record39_rec_valid <= 1'd0;
		main_rtio_core_outputs_record40_rec_valid <= 1'd0;
		main_rtio_core_outputs_record41_rec_valid <= 1'd0;
		main_rtio_core_outputs_record42_rec_valid <= 1'd0;
		main_rtio_core_outputs_record43_rec_valid <= 1'd0;
		main_rtio_core_outputs_record44_rec_valid <= 1'd0;
		main_rtio_core_outputs_record45_rec_valid <= 1'd0;
		main_rtio_core_outputs_record46_rec_valid <= 1'd0;
		main_rtio_core_outputs_record47_rec_valid <= 1'd0;
		main_rtio_core_outputs_record0_valid1 <= 1'd0;
		main_rtio_core_outputs_record1_valid1 <= 1'd0;
		main_rtio_core_outputs_record2_valid1 <= 1'd0;
		main_rtio_core_outputs_record3_valid1 <= 1'd0;
		main_rtio_core_outputs_record4_valid1 <= 1'd0;
		main_rtio_core_outputs_record5_valid1 <= 1'd0;
		main_rtio_core_outputs_record6_valid1 <= 1'd0;
		main_rtio_core_outputs_record7_valid1 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r0 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r0 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r1 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r1 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r2 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r2 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r3 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r3 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r4 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r4 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r5 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r5 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r6 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r6 <= 1'd0;
		main_rtio_core_outputs_replace_occured_r7 <= 1'd0;
		main_rtio_core_outputs_nondata_replace_occured_r7 <= 1'd0;
		main_rtio_core_outputs_stb_r0 <= 1'd0;
		main_rtio_core_outputs_stb_r1 <= 1'd0;
		main_rtio_core_outputs_stb_r2 <= 1'd0;
		main_rtio_core_outputs_stb_r3 <= 1'd0;
		main_rtio_core_outputs_stb_r4 <= 1'd0;
		main_rtio_core_outputs_stb_r5 <= 1'd0;
		main_rtio_core_outputs_stb_r6 <= 1'd0;
		main_rtio_core_outputs_stb_r7 <= 1'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter0_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter0_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer0_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter2_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter2_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer1_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter4_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter4_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer2_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter6_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter6_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer3_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter8_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter8_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer4_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter10_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter10_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer5_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter12_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter12_q_binary <= 10'd0;
		main_rtio_core_inputs_blindtransfer6_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter14_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter14_q_binary <= 3'd0;
		main_rtio_core_inputs_blindtransfer7_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter16_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter16_q_binary <= 8'd0;
		main_rtio_core_inputs_blindtransfer8_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter18_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter18_q_binary <= 8'd0;
		main_rtio_core_inputs_blindtransfer9_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter20_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter20_q_binary <= 8'd0;
		main_rtio_core_inputs_blindtransfer10_blind <= 1'd0;
		main_rtio_core_inputs_asyncfifo11_graycounter22_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo11_graycounter22_q_binary <= 3'd0;
		main_rtio_core_inputs_blindtransfer11_blind <= 1'd0;
		main_rtio_core_o_collision_sync_blind <= 1'd0;
		main_rtio_core_o_busy_sync_blind <= 1'd0;
		main_mon_bussynchronizer28_starter <= 1'd1;
		main_mon_bussynchronizer28_count <= 8'd128;
		main_mon_bussynchronizer29_starter <= 1'd1;
		main_mon_bussynchronizer29_count <= 8'd128;
		main_mon_bussynchronizer30_starter <= 1'd1;
		main_mon_bussynchronizer30_count <= 8'd128;
		main_mon_bussynchronizer31_starter <= 1'd1;
		main_mon_bussynchronizer31_count <= 8'd128;
		main_mon_bussynchronizer32_starter <= 1'd1;
		main_mon_bussynchronizer32_count <= 8'd128;
		main_mon_bussynchronizer33_starter <= 1'd1;
		main_mon_bussynchronizer33_count <= 8'd128;
		main_mon_bussynchronizer34_starter <= 1'd1;
		main_mon_bussynchronizer34_count <= 8'd128;
		main_mon_bussynchronizer35_starter <= 1'd1;
		main_mon_bussynchronizer35_count <= 8'd128;
		main_mon_bussynchronizer36_starter <= 1'd1;
		main_mon_bussynchronizer36_count <= 8'd128;
		main_mon_bussynchronizer37_starter <= 1'd1;
		main_mon_bussynchronizer37_count <= 8'd128;
		main_mon_bussynchronizer38_starter <= 1'd1;
		main_mon_bussynchronizer38_count <= 8'd128;
	end
	builder_xilinxmultiregimpl12_regs0 <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q;
	builder_xilinxmultiregimpl12_regs1 <= builder_xilinxmultiregimpl12_regs0;
	builder_xilinxmultiregimpl14_regs0 <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q;
	builder_xilinxmultiregimpl14_regs1 <= builder_xilinxmultiregimpl14_regs0;
	builder_xilinxmultiregimpl16_regs0 <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q;
	builder_xilinxmultiregimpl16_regs1 <= builder_xilinxmultiregimpl16_regs0;
	builder_xilinxmultiregimpl18_regs0 <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q;
	builder_xilinxmultiregimpl18_regs1 <= builder_xilinxmultiregimpl18_regs0;
	builder_xilinxmultiregimpl20_regs0 <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q;
	builder_xilinxmultiregimpl20_regs1 <= builder_xilinxmultiregimpl20_regs0;
	builder_xilinxmultiregimpl22_regs0 <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q;
	builder_xilinxmultiregimpl22_regs1 <= builder_xilinxmultiregimpl22_regs0;
	builder_xilinxmultiregimpl24_regs0 <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q;
	builder_xilinxmultiregimpl24_regs1 <= builder_xilinxmultiregimpl24_regs0;
	builder_xilinxmultiregimpl26_regs0 <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q;
	builder_xilinxmultiregimpl26_regs1 <= builder_xilinxmultiregimpl26_regs0;
	builder_xilinxmultiregimpl29_regs0 <= main_rtio_core_inputs_asyncfifo0_graycounter1_q;
	builder_xilinxmultiregimpl29_regs1 <= builder_xilinxmultiregimpl29_regs0;
	builder_xilinxmultiregimpl31_regs0 <= main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i;
	builder_xilinxmultiregimpl31_regs1 <= builder_xilinxmultiregimpl31_regs0;
	builder_xilinxmultiregimpl33_regs0 <= main_rtio_core_inputs_asyncfifo1_graycounter3_q;
	builder_xilinxmultiregimpl33_regs1 <= builder_xilinxmultiregimpl33_regs0;
	builder_xilinxmultiregimpl35_regs0 <= main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i;
	builder_xilinxmultiregimpl35_regs1 <= builder_xilinxmultiregimpl35_regs0;
	builder_xilinxmultiregimpl37_regs0 <= main_rtio_core_inputs_asyncfifo2_graycounter5_q;
	builder_xilinxmultiregimpl37_regs1 <= builder_xilinxmultiregimpl37_regs0;
	builder_xilinxmultiregimpl39_regs0 <= main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i;
	builder_xilinxmultiregimpl39_regs1 <= builder_xilinxmultiregimpl39_regs0;
	builder_xilinxmultiregimpl41_regs0 <= main_rtio_core_inputs_asyncfifo3_graycounter7_q;
	builder_xilinxmultiregimpl41_regs1 <= builder_xilinxmultiregimpl41_regs0;
	builder_xilinxmultiregimpl43_regs0 <= main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i;
	builder_xilinxmultiregimpl43_regs1 <= builder_xilinxmultiregimpl43_regs0;
	builder_xilinxmultiregimpl45_regs0 <= main_rtio_core_inputs_asyncfifo4_graycounter9_q;
	builder_xilinxmultiregimpl45_regs1 <= builder_xilinxmultiregimpl45_regs0;
	builder_xilinxmultiregimpl47_regs0 <= main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i;
	builder_xilinxmultiregimpl47_regs1 <= builder_xilinxmultiregimpl47_regs0;
	builder_xilinxmultiregimpl49_regs0 <= main_rtio_core_inputs_asyncfifo5_graycounter11_q;
	builder_xilinxmultiregimpl49_regs1 <= builder_xilinxmultiregimpl49_regs0;
	builder_xilinxmultiregimpl51_regs0 <= main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i;
	builder_xilinxmultiregimpl51_regs1 <= builder_xilinxmultiregimpl51_regs0;
	builder_xilinxmultiregimpl53_regs0 <= main_rtio_core_inputs_asyncfifo6_graycounter13_q;
	builder_xilinxmultiregimpl53_regs1 <= builder_xilinxmultiregimpl53_regs0;
	builder_xilinxmultiregimpl55_regs0 <= main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i;
	builder_xilinxmultiregimpl55_regs1 <= builder_xilinxmultiregimpl55_regs0;
	builder_xilinxmultiregimpl57_regs0 <= main_rtio_core_inputs_asyncfifo7_graycounter15_q;
	builder_xilinxmultiregimpl57_regs1 <= builder_xilinxmultiregimpl57_regs0;
	builder_xilinxmultiregimpl59_regs0 <= main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i;
	builder_xilinxmultiregimpl59_regs1 <= builder_xilinxmultiregimpl59_regs0;
	builder_xilinxmultiregimpl61_regs0 <= main_rtio_core_inputs_asyncfifo8_graycounter17_q;
	builder_xilinxmultiregimpl61_regs1 <= builder_xilinxmultiregimpl61_regs0;
	builder_xilinxmultiregimpl63_regs0 <= main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i;
	builder_xilinxmultiregimpl63_regs1 <= builder_xilinxmultiregimpl63_regs0;
	builder_xilinxmultiregimpl65_regs0 <= main_rtio_core_inputs_asyncfifo9_graycounter19_q;
	builder_xilinxmultiregimpl65_regs1 <= builder_xilinxmultiregimpl65_regs0;
	builder_xilinxmultiregimpl67_regs0 <= main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i;
	builder_xilinxmultiregimpl67_regs1 <= builder_xilinxmultiregimpl67_regs0;
	builder_xilinxmultiregimpl69_regs0 <= main_rtio_core_inputs_asyncfifo10_graycounter21_q;
	builder_xilinxmultiregimpl69_regs1 <= builder_xilinxmultiregimpl69_regs0;
	builder_xilinxmultiregimpl71_regs0 <= main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i;
	builder_xilinxmultiregimpl71_regs1 <= builder_xilinxmultiregimpl71_regs0;
	builder_xilinxmultiregimpl73_regs0 <= main_rtio_core_inputs_asyncfifo11_graycounter23_q;
	builder_xilinxmultiregimpl73_regs1 <= builder_xilinxmultiregimpl73_regs0;
	builder_xilinxmultiregimpl75_regs0 <= main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_i;
	builder_xilinxmultiregimpl75_regs1 <= builder_xilinxmultiregimpl75_regs0;
	builder_xilinxmultiregimpl77_regs0 <= main_rtio_core_o_collision_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl77_regs1 <= builder_xilinxmultiregimpl77_regs0;
	builder_xilinxmultiregimpl80_regs0 <= main_rtio_core_o_busy_sync_ps_ack_toggle_i;
	builder_xilinxmultiregimpl80_regs1 <= builder_xilinxmultiregimpl80_regs0;
	builder_xilinxmultiregimpl111_regs0 <= main_mon_bussynchronizer28_pong_toggle_i;
	builder_xilinxmultiregimpl111_regs1 <= builder_xilinxmultiregimpl111_regs0;
	builder_xilinxmultiregimpl114_regs0 <= main_mon_bussynchronizer29_pong_toggle_i;
	builder_xilinxmultiregimpl114_regs1 <= builder_xilinxmultiregimpl114_regs0;
	builder_xilinxmultiregimpl117_regs0 <= main_mon_bussynchronizer30_pong_toggle_i;
	builder_xilinxmultiregimpl117_regs1 <= builder_xilinxmultiregimpl117_regs0;
	builder_xilinxmultiregimpl120_regs0 <= main_mon_bussynchronizer31_pong_toggle_i;
	builder_xilinxmultiregimpl120_regs1 <= builder_xilinxmultiregimpl120_regs0;
	builder_xilinxmultiregimpl123_regs0 <= main_mon_bussynchronizer32_pong_toggle_i;
	builder_xilinxmultiregimpl123_regs1 <= builder_xilinxmultiregimpl123_regs0;
	builder_xilinxmultiregimpl126_regs0 <= main_mon_bussynchronizer33_pong_toggle_i;
	builder_xilinxmultiregimpl126_regs1 <= builder_xilinxmultiregimpl126_regs0;
	builder_xilinxmultiregimpl129_regs0 <= main_mon_bussynchronizer34_pong_toggle_i;
	builder_xilinxmultiregimpl129_regs1 <= builder_xilinxmultiregimpl129_regs0;
	builder_xilinxmultiregimpl132_regs0 <= main_mon_bussynchronizer35_pong_toggle_i;
	builder_xilinxmultiregimpl132_regs1 <= builder_xilinxmultiregimpl132_regs0;
	builder_xilinxmultiregimpl135_regs0 <= main_mon_bussynchronizer36_pong_toggle_i;
	builder_xilinxmultiregimpl135_regs1 <= builder_xilinxmultiregimpl135_regs0;
	builder_xilinxmultiregimpl138_regs0 <= main_mon_bussynchronizer37_pong_toggle_i;
	builder_xilinxmultiregimpl138_regs1 <= builder_xilinxmultiregimpl138_regs0;
	builder_xilinxmultiregimpl141_regs0 <= main_mon_bussynchronizer38_pong_toggle_i;
	builder_xilinxmultiregimpl141_regs1 <= builder_xilinxmultiregimpl141_regs0;
	builder_xilinxmultiregimpl143_regs0 <= main_inj_o_sys0;
	builder_xilinxmultiregimpl143_regs1 <= builder_xilinxmultiregimpl143_regs0;
	builder_xilinxmultiregimpl144_regs0 <= main_inj_o_sys1;
	builder_xilinxmultiregimpl144_regs1 <= builder_xilinxmultiregimpl144_regs0;
	builder_xilinxmultiregimpl145_regs0 <= main_inj_o_sys2;
	builder_xilinxmultiregimpl145_regs1 <= builder_xilinxmultiregimpl145_regs0;
	builder_xilinxmultiregimpl146_regs0 <= main_inj_o_sys3;
	builder_xilinxmultiregimpl146_regs1 <= builder_xilinxmultiregimpl146_regs0;
	builder_xilinxmultiregimpl147_regs0 <= main_inj_o_sys4;
	builder_xilinxmultiregimpl147_regs1 <= builder_xilinxmultiregimpl147_regs0;
	builder_xilinxmultiregimpl148_regs0 <= main_inj_o_sys5;
	builder_xilinxmultiregimpl148_regs1 <= builder_xilinxmultiregimpl148_regs0;
	builder_xilinxmultiregimpl149_regs0 <= main_inj_o_sys6;
	builder_xilinxmultiregimpl149_regs1 <= builder_xilinxmultiregimpl149_regs0;
	builder_xilinxmultiregimpl150_regs0 <= main_inj_o_sys7;
	builder_xilinxmultiregimpl150_regs1 <= builder_xilinxmultiregimpl150_regs0;
	builder_xilinxmultiregimpl151_regs0 <= main_inj_o_sys8;
	builder_xilinxmultiregimpl151_regs1 <= builder_xilinxmultiregimpl151_regs0;
	builder_xilinxmultiregimpl152_regs0 <= main_inj_o_sys9;
	builder_xilinxmultiregimpl152_regs1 <= builder_xilinxmultiregimpl152_regs0;
	builder_xilinxmultiregimpl153_regs0 <= main_inj_o_sys10;
	builder_xilinxmultiregimpl153_regs1 <= builder_xilinxmultiregimpl153_regs0;
	builder_xilinxmultiregimpl154_regs0 <= main_inj_o_sys11;
	builder_xilinxmultiregimpl154_regs1 <= builder_xilinxmultiregimpl154_regs0;
	builder_xilinxmultiregimpl155_regs0 <= main_inj_o_sys12;
	builder_xilinxmultiregimpl155_regs1 <= builder_xilinxmultiregimpl155_regs0;
	builder_xilinxmultiregimpl156_regs0 <= main_inj_o_sys13;
	builder_xilinxmultiregimpl156_regs1 <= builder_xilinxmultiregimpl156_regs0;
	builder_xilinxmultiregimpl157_regs0 <= main_inj_o_sys14;
	builder_xilinxmultiregimpl157_regs1 <= builder_xilinxmultiregimpl157_regs0;
	builder_xilinxmultiregimpl158_regs0 <= main_inj_o_sys15;
	builder_xilinxmultiregimpl158_regs1 <= builder_xilinxmultiregimpl158_regs0;
	builder_xilinxmultiregimpl159_regs0 <= main_inj_o_sys16;
	builder_xilinxmultiregimpl159_regs1 <= builder_xilinxmultiregimpl159_regs0;
	builder_xilinxmultiregimpl160_regs0 <= main_inj_o_sys17;
	builder_xilinxmultiregimpl160_regs1 <= builder_xilinxmultiregimpl160_regs0;
	builder_xilinxmultiregimpl161_regs0 <= main_inj_o_sys18;
	builder_xilinxmultiregimpl161_regs1 <= builder_xilinxmultiregimpl161_regs0;
	builder_xilinxmultiregimpl162_regs0 <= main_inj_o_sys19;
	builder_xilinxmultiregimpl162_regs1 <= builder_xilinxmultiregimpl162_regs0;
	builder_xilinxmultiregimpl163_regs0 <= main_inj_o_sys20;
	builder_xilinxmultiregimpl163_regs1 <= builder_xilinxmultiregimpl163_regs0;
	builder_xilinxmultiregimpl164_regs0 <= main_inj_o_sys21;
	builder_xilinxmultiregimpl164_regs1 <= builder_xilinxmultiregimpl164_regs0;
	builder_xilinxmultiregimpl165_regs0 <= main_inj_o_sys22;
	builder_xilinxmultiregimpl165_regs1 <= builder_xilinxmultiregimpl165_regs0;
	builder_xilinxmultiregimpl166_regs0 <= main_inj_o_sys23;
	builder_xilinxmultiregimpl166_regs1 <= builder_xilinxmultiregimpl166_regs0;
	builder_xilinxmultiregimpl167_regs0 <= main_inj_o_sys24;
	builder_xilinxmultiregimpl167_regs1 <= builder_xilinxmultiregimpl167_regs0;
	builder_xilinxmultiregimpl168_regs0 <= main_inj_o_sys25;
	builder_xilinxmultiregimpl168_regs1 <= builder_xilinxmultiregimpl168_regs0;
	builder_xilinxmultiregimpl169_regs0 <= main_inj_o_sys26;
	builder_xilinxmultiregimpl169_regs1 <= builder_xilinxmultiregimpl169_regs0;
	builder_xilinxmultiregimpl170_regs0 <= main_inj_o_sys27;
	builder_xilinxmultiregimpl170_regs1 <= builder_xilinxmultiregimpl170_regs0;
	builder_xilinxmultiregimpl171_regs0 <= main_inj_o_sys28;
	builder_xilinxmultiregimpl171_regs1 <= builder_xilinxmultiregimpl171_regs0;
	builder_xilinxmultiregimpl172_regs0 <= main_inj_o_sys29;
	builder_xilinxmultiregimpl172_regs1 <= builder_xilinxmultiregimpl172_regs0;
	builder_xilinxmultiregimpl173_regs0 <= main_inj_o_sys30;
	builder_xilinxmultiregimpl173_regs1 <= builder_xilinxmultiregimpl173_regs0;
	builder_xilinxmultiregimpl174_regs0 <= main_inj_o_sys31;
	builder_xilinxmultiregimpl174_regs1 <= builder_xilinxmultiregimpl174_regs0;
	builder_xilinxmultiregimpl175_regs0 <= main_inj_o_sys32;
	builder_xilinxmultiregimpl175_regs1 <= builder_xilinxmultiregimpl175_regs0;
	builder_xilinxmultiregimpl176_regs0 <= main_inj_o_sys33;
	builder_xilinxmultiregimpl176_regs1 <= builder_xilinxmultiregimpl176_regs0;
	builder_xilinxmultiregimpl177_regs0 <= main_inj_o_sys34;
	builder_xilinxmultiregimpl177_regs1 <= builder_xilinxmultiregimpl177_regs0;
	builder_xilinxmultiregimpl178_regs0 <= main_inj_o_sys35;
	builder_xilinxmultiregimpl178_regs1 <= builder_xilinxmultiregimpl178_regs0;
	builder_xilinxmultiregimpl179_regs0 <= main_inj_o_sys36;
	builder_xilinxmultiregimpl179_regs1 <= builder_xilinxmultiregimpl179_regs0;
	builder_xilinxmultiregimpl180_regs0 <= main_inj_o_sys37;
	builder_xilinxmultiregimpl180_regs1 <= builder_xilinxmultiregimpl180_regs0;
	builder_xilinxmultiregimpl181_regs0 <= main_inj_o_sys38;
	builder_xilinxmultiregimpl181_regs1 <= builder_xilinxmultiregimpl181_regs0;
	builder_xilinxmultiregimpl182_regs0 <= main_inj_o_sys39;
	builder_xilinxmultiregimpl182_regs1 <= builder_xilinxmultiregimpl182_regs0;
	builder_xilinxmultiregimpl183_regs0 <= main_inj_o_sys40;
	builder_xilinxmultiregimpl183_regs1 <= builder_xilinxmultiregimpl183_regs0;
	builder_xilinxmultiregimpl184_regs0 <= main_inj_o_sys41;
	builder_xilinxmultiregimpl184_regs1 <= builder_xilinxmultiregimpl184_regs0;
	builder_xilinxmultiregimpl185_regs0 <= main_inj_o_sys42;
	builder_xilinxmultiregimpl185_regs1 <= builder_xilinxmultiregimpl185_regs0;
	builder_xilinxmultiregimpl186_regs0 <= main_inj_o_sys43;
	builder_xilinxmultiregimpl186_regs1 <= builder_xilinxmultiregimpl186_regs0;
	builder_xilinxmultiregimpl187_regs0 <= main_inj_o_sys44;
	builder_xilinxmultiregimpl187_regs1 <= builder_xilinxmultiregimpl187_regs0;
	builder_xilinxmultiregimpl188_regs0 <= main_inj_o_sys45;
	builder_xilinxmultiregimpl188_regs1 <= builder_xilinxmultiregimpl188_regs0;
	builder_xilinxmultiregimpl189_regs0 <= main_inj_o_sys46;
	builder_xilinxmultiregimpl189_regs1 <= builder_xilinxmultiregimpl189_regs0;
	builder_xilinxmultiregimpl190_regs0 <= main_inj_o_sys47;
	builder_xilinxmultiregimpl190_regs1 <= builder_xilinxmultiregimpl190_regs0;
	builder_xilinxmultiregimpl191_regs0 <= main_inj_o_sys48;
	builder_xilinxmultiregimpl191_regs1 <= builder_xilinxmultiregimpl191_regs0;
end

always @(posedge rio_phy_clk) begin
	if (main_output_8x0_stb) begin
		main_output_8x0_previous_data <= main_output_8x0_data;
	end
	if (main_output_8x0_override_en) begin
		main_output_8x0_o <= {8{main_output_8x0_override_o}};
	end else begin
		if (((main_output_8x0_stb & (~main_output_8x0_previous_data)) & main_output_8x0_data)) begin
			main_output_8x0_o <= builder_sync_f_t_array_muxed0;
		end else begin
			if (((main_output_8x0_stb & main_output_8x0_previous_data) & (~main_output_8x0_data))) begin
				main_output_8x0_o <= builder_sync_f_f_array_muxed0;
			end else begin
				main_output_8x0_o <= {8{main_output_8x0_previous_data}};
			end
		end
	end
	if (main_output_8x1_stb) begin
		main_output_8x1_previous_data <= main_output_8x1_data;
	end
	if (main_output_8x1_override_en) begin
		main_output_8x1_o <= {8{main_output_8x1_override_o}};
	end else begin
		if (((main_output_8x1_stb & (~main_output_8x1_previous_data)) & main_output_8x1_data)) begin
			main_output_8x1_o <= builder_sync_f_t_array_muxed1;
		end else begin
			if (((main_output_8x1_stb & main_output_8x1_previous_data) & (~main_output_8x1_data))) begin
				main_output_8x1_o <= builder_sync_f_f_array_muxed1;
			end else begin
				main_output_8x1_o <= {8{main_output_8x1_previous_data}};
			end
		end
	end
	if (main_output_8x2_stb) begin
		main_output_8x2_previous_data <= main_output_8x2_data;
	end
	if (main_output_8x2_override_en) begin
		main_output_8x2_o <= {8{main_output_8x2_override_o}};
	end else begin
		if (((main_output_8x2_stb & (~main_output_8x2_previous_data)) & main_output_8x2_data)) begin
			main_output_8x2_o <= builder_sync_f_t_array_muxed2;
		end else begin
			if (((main_output_8x2_stb & main_output_8x2_previous_data) & (~main_output_8x2_data))) begin
				main_output_8x2_o <= builder_sync_f_f_array_muxed2;
			end else begin
				main_output_8x2_o <= {8{main_output_8x2_previous_data}};
			end
		end
	end
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd1))) begin
		main_inout_8x0_inout_8x0_oe_k <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_inout_8x0_oe <= main_inout_8x0_inout_8x0_override_oe;
	end else begin
		main_inout_8x0_inout_8x0_oe <= main_inout_8x0_inout_8x0_oe_k;
	end
	main_inout_8x0_inout_8x0_i_d <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_stb <= ((main_inout_8x0_inout_8x0_sample | (main_inout_8x0_inout_8x0_sensitivity[0] & (main_inout_8x0_serdes_i0[7] & (~main_inout_8x0_inout_8x0_i_d)))) | (main_inout_8x0_inout_8x0_sensitivity[1] & ((~main_inout_8x0_serdes_i0[7]) & main_inout_8x0_inout_8x0_i_d)));
	main_inout_8x0_inout_8x0_iinterface0_data <= main_inout_8x0_serdes_i0[7];
	main_inout_8x0_inout_8x0_iinterface0_fine_ts <= main_inout_8x0_inout_8x0_o;
	if ((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0))) begin
		main_inout_8x0_inout_8x0_previous_data <= main_inout_8x0_inout_8x0_ointerface0_data[0];
	end
	if (main_inout_8x0_inout_8x0_override_en) begin
		main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_override_o}};
	end else begin
		if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & (~main_inout_8x0_inout_8x0_previous_data)) & main_inout_8x0_inout_8x0_ointerface0_data[0])) begin
			main_inout_8x0_serdes_o0 <= builder_sync_f_t_array_muxed3;
		end else begin
			if ((((main_inout_8x0_inout_8x0_ointerface0_stb & (main_inout_8x0_inout_8x0_ointerface0_address == 1'd0)) & main_inout_8x0_inout_8x0_previous_data) & (~main_inout_8x0_inout_8x0_ointerface0_data[0]))) begin
				main_inout_8x0_serdes_o0 <= builder_sync_f_f_array_muxed3;
			end else begin
				main_inout_8x0_serdes_o0 <= {8{main_inout_8x0_inout_8x0_previous_data}};
			end
		end
	end
	if (main_output_8x3_stb) begin
		main_output_8x3_previous_data <= main_output_8x3_data;
	end
	if (main_output_8x3_override_en) begin
		main_output_8x3_o <= {8{main_output_8x3_override_o}};
	end else begin
		if (((main_output_8x3_stb & (~main_output_8x3_previous_data)) & main_output_8x3_data)) begin
			main_output_8x3_o <= builder_sync_f_t_array_muxed4;
		end else begin
			if (((main_output_8x3_stb & main_output_8x3_previous_data) & (~main_output_8x3_data))) begin
				main_output_8x3_o <= builder_sync_f_f_array_muxed4;
			end else begin
				main_output_8x3_o <= {8{main_output_8x3_previous_data}};
			end
		end
	end
	if (main_output_8x4_stb) begin
		main_output_8x4_previous_data <= main_output_8x4_data;
	end
	if (main_output_8x4_override_en) begin
		main_output_8x4_o <= {8{main_output_8x4_override_o}};
	end else begin
		if (((main_output_8x4_stb & (~main_output_8x4_previous_data)) & main_output_8x4_data)) begin
			main_output_8x4_o <= builder_sync_f_t_array_muxed5;
		end else begin
			if (((main_output_8x4_stb & main_output_8x4_previous_data) & (~main_output_8x4_data))) begin
				main_output_8x4_o <= builder_sync_f_f_array_muxed5;
			end else begin
				main_output_8x4_o <= {8{main_output_8x4_previous_data}};
			end
		end
	end
	if (main_output_8x5_stb) begin
		main_output_8x5_previous_data <= main_output_8x5_data;
	end
	if (main_output_8x5_override_en) begin
		main_output_8x5_o <= {8{main_output_8x5_override_o}};
	end else begin
		if (((main_output_8x5_stb & (~main_output_8x5_previous_data)) & main_output_8x5_data)) begin
			main_output_8x5_o <= builder_sync_f_t_array_muxed6;
		end else begin
			if (((main_output_8x5_stb & main_output_8x5_previous_data) & (~main_output_8x5_data))) begin
				main_output_8x5_o <= builder_sync_f_f_array_muxed6;
			end else begin
				main_output_8x5_o <= {8{main_output_8x5_previous_data}};
			end
		end
	end
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd1))) begin
		main_inout_8x1_inout_8x1_oe_k <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_inout_8x1_oe <= main_inout_8x1_inout_8x1_override_oe;
	end else begin
		main_inout_8x1_inout_8x1_oe <= main_inout_8x1_inout_8x1_oe_k;
	end
	main_inout_8x1_inout_8x1_i_d <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_stb <= ((main_inout_8x1_inout_8x1_sample | (main_inout_8x1_inout_8x1_sensitivity[0] & (main_inout_8x1_serdes_i0[7] & (~main_inout_8x1_inout_8x1_i_d)))) | (main_inout_8x1_inout_8x1_sensitivity[1] & ((~main_inout_8x1_serdes_i0[7]) & main_inout_8x1_inout_8x1_i_d)));
	main_inout_8x1_inout_8x1_iinterface1_data <= main_inout_8x1_serdes_i0[7];
	main_inout_8x1_inout_8x1_iinterface1_fine_ts <= main_inout_8x1_inout_8x1_o;
	if ((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0))) begin
		main_inout_8x1_inout_8x1_previous_data <= main_inout_8x1_inout_8x1_ointerface1_data[0];
	end
	if (main_inout_8x1_inout_8x1_override_en) begin
		main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_override_o}};
	end else begin
		if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & (~main_inout_8x1_inout_8x1_previous_data)) & main_inout_8x1_inout_8x1_ointerface1_data[0])) begin
			main_inout_8x1_serdes_o0 <= builder_sync_f_t_array_muxed7;
		end else begin
			if ((((main_inout_8x1_inout_8x1_ointerface1_stb & (main_inout_8x1_inout_8x1_ointerface1_address == 1'd0)) & main_inout_8x1_inout_8x1_previous_data) & (~main_inout_8x1_inout_8x1_ointerface1_data[0]))) begin
				main_inout_8x1_serdes_o0 <= builder_sync_f_f_array_muxed7;
			end else begin
				main_inout_8x1_serdes_o0 <= {8{main_inout_8x1_inout_8x1_previous_data}};
			end
		end
	end
	if (main_output_8x6_stb) begin
		main_output_8x6_previous_data <= main_output_8x6_data;
	end
	if (main_output_8x6_override_en) begin
		main_output_8x6_o <= {8{main_output_8x6_override_o}};
	end else begin
		if (((main_output_8x6_stb & (~main_output_8x6_previous_data)) & main_output_8x6_data)) begin
			main_output_8x6_o <= builder_sync_f_t_array_muxed8;
		end else begin
			if (((main_output_8x6_stb & main_output_8x6_previous_data) & (~main_output_8x6_data))) begin
				main_output_8x6_o <= builder_sync_f_f_array_muxed8;
			end else begin
				main_output_8x6_o <= {8{main_output_8x6_previous_data}};
			end
		end
	end
	if (main_output_8x7_stb) begin
		main_output_8x7_previous_data <= main_output_8x7_data;
	end
	if (main_output_8x7_override_en) begin
		main_output_8x7_o <= {8{main_output_8x7_override_o}};
	end else begin
		if (((main_output_8x7_stb & (~main_output_8x7_previous_data)) & main_output_8x7_data)) begin
			main_output_8x7_o <= builder_sync_f_t_array_muxed9;
		end else begin
			if (((main_output_8x7_stb & main_output_8x7_previous_data) & (~main_output_8x7_data))) begin
				main_output_8x7_o <= builder_sync_f_f_array_muxed9;
			end else begin
				main_output_8x7_o <= {8{main_output_8x7_previous_data}};
			end
		end
	end
	if (main_output_8x8_stb) begin
		main_output_8x8_previous_data <= main_output_8x8_data;
	end
	if (main_output_8x8_override_en) begin
		main_output_8x8_o <= {8{main_output_8x8_override_o}};
	end else begin
		if (((main_output_8x8_stb & (~main_output_8x8_previous_data)) & main_output_8x8_data)) begin
			main_output_8x8_o <= builder_sync_f_t_array_muxed10;
		end else begin
			if (((main_output_8x8_stb & main_output_8x8_previous_data) & (~main_output_8x8_data))) begin
				main_output_8x8_o <= builder_sync_f_f_array_muxed10;
			end else begin
				main_output_8x8_o <= {8{main_output_8x8_previous_data}};
			end
		end
	end
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd1))) begin
		main_inout_8x2_inout_8x2_oe_k <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_inout_8x2_oe <= main_inout_8x2_inout_8x2_override_oe;
	end else begin
		main_inout_8x2_inout_8x2_oe <= main_inout_8x2_inout_8x2_oe_k;
	end
	main_inout_8x2_inout_8x2_i_d <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_stb <= ((main_inout_8x2_inout_8x2_sample | (main_inout_8x2_inout_8x2_sensitivity[0] & (main_inout_8x2_serdes_i0[7] & (~main_inout_8x2_inout_8x2_i_d)))) | (main_inout_8x2_inout_8x2_sensitivity[1] & ((~main_inout_8x2_serdes_i0[7]) & main_inout_8x2_inout_8x2_i_d)));
	main_inout_8x2_inout_8x2_iinterface2_data <= main_inout_8x2_serdes_i0[7];
	main_inout_8x2_inout_8x2_iinterface2_fine_ts <= main_inout_8x2_inout_8x2_o;
	if ((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0))) begin
		main_inout_8x2_inout_8x2_previous_data <= main_inout_8x2_inout_8x2_ointerface2_data[0];
	end
	if (main_inout_8x2_inout_8x2_override_en) begin
		main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_override_o}};
	end else begin
		if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & (~main_inout_8x2_inout_8x2_previous_data)) & main_inout_8x2_inout_8x2_ointerface2_data[0])) begin
			main_inout_8x2_serdes_o0 <= builder_sync_f_t_array_muxed11;
		end else begin
			if ((((main_inout_8x2_inout_8x2_ointerface2_stb & (main_inout_8x2_inout_8x2_ointerface2_address == 1'd0)) & main_inout_8x2_inout_8x2_previous_data) & (~main_inout_8x2_inout_8x2_ointerface2_data[0]))) begin
				main_inout_8x2_serdes_o0 <= builder_sync_f_f_array_muxed11;
			end else begin
				main_inout_8x2_serdes_o0 <= {8{main_inout_8x2_inout_8x2_previous_data}};
			end
		end
	end
	if (main_output_8x9_stb) begin
		main_output_8x9_previous_data <= main_output_8x9_data;
	end
	if (main_output_8x9_override_en) begin
		main_output_8x9_o <= {8{main_output_8x9_override_o}};
	end else begin
		if (((main_output_8x9_stb & (~main_output_8x9_previous_data)) & main_output_8x9_data)) begin
			main_output_8x9_o <= builder_sync_f_t_array_muxed12;
		end else begin
			if (((main_output_8x9_stb & main_output_8x9_previous_data) & (~main_output_8x9_data))) begin
				main_output_8x9_o <= builder_sync_f_f_array_muxed12;
			end else begin
				main_output_8x9_o <= {8{main_output_8x9_previous_data}};
			end
		end
	end
	if (main_output_8x10_stb) begin
		main_output_8x10_previous_data <= main_output_8x10_data;
	end
	if (main_output_8x10_override_en) begin
		main_output_8x10_o <= {8{main_output_8x10_override_o}};
	end else begin
		if (((main_output_8x10_stb & (~main_output_8x10_previous_data)) & main_output_8x10_data)) begin
			main_output_8x10_o <= builder_sync_f_t_array_muxed13;
		end else begin
			if (((main_output_8x10_stb & main_output_8x10_previous_data) & (~main_output_8x10_data))) begin
				main_output_8x10_o <= builder_sync_f_f_array_muxed13;
			end else begin
				main_output_8x10_o <= {8{main_output_8x10_previous_data}};
			end
		end
	end
	if (main_output_8x11_stb) begin
		main_output_8x11_previous_data <= main_output_8x11_data;
	end
	if (main_output_8x11_override_en) begin
		main_output_8x11_o <= {8{main_output_8x11_override_o}};
	end else begin
		if (((main_output_8x11_stb & (~main_output_8x11_previous_data)) & main_output_8x11_data)) begin
			main_output_8x11_o <= builder_sync_f_t_array_muxed14;
		end else begin
			if (((main_output_8x11_stb & main_output_8x11_previous_data) & (~main_output_8x11_data))) begin
				main_output_8x11_o <= builder_sync_f_f_array_muxed14;
			end else begin
				main_output_8x11_o <= {8{main_output_8x11_previous_data}};
			end
		end
	end
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd1))) begin
		main_inout_8x3_inout_8x3_oe_k <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_inout_8x3_oe <= main_inout_8x3_inout_8x3_override_oe;
	end else begin
		main_inout_8x3_inout_8x3_oe <= main_inout_8x3_inout_8x3_oe_k;
	end
	main_inout_8x3_inout_8x3_i_d <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_stb <= ((main_inout_8x3_inout_8x3_sample | (main_inout_8x3_inout_8x3_sensitivity[0] & (main_inout_8x3_serdes_i0[7] & (~main_inout_8x3_inout_8x3_i_d)))) | (main_inout_8x3_inout_8x3_sensitivity[1] & ((~main_inout_8x3_serdes_i0[7]) & main_inout_8x3_inout_8x3_i_d)));
	main_inout_8x3_inout_8x3_iinterface3_data <= main_inout_8x3_serdes_i0[7];
	main_inout_8x3_inout_8x3_iinterface3_fine_ts <= main_inout_8x3_inout_8x3_o;
	if ((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0))) begin
		main_inout_8x3_inout_8x3_previous_data <= main_inout_8x3_inout_8x3_ointerface3_data[0];
	end
	if (main_inout_8x3_inout_8x3_override_en) begin
		main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_override_o}};
	end else begin
		if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & (~main_inout_8x3_inout_8x3_previous_data)) & main_inout_8x3_inout_8x3_ointerface3_data[0])) begin
			main_inout_8x3_serdes_o0 <= builder_sync_f_t_array_muxed15;
		end else begin
			if ((((main_inout_8x3_inout_8x3_ointerface3_stb & (main_inout_8x3_inout_8x3_ointerface3_address == 1'd0)) & main_inout_8x3_inout_8x3_previous_data) & (~main_inout_8x3_inout_8x3_ointerface3_data[0]))) begin
				main_inout_8x3_serdes_o0 <= builder_sync_f_f_array_muxed15;
			end else begin
				main_inout_8x3_serdes_o0 <= {8{main_inout_8x3_inout_8x3_previous_data}};
			end
		end
	end
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd1))) begin
		main_inout_8x4_inout_8x4_oe_k <= main_inout_8x4_inout_8x4_ointerface4_data[0];
	end
	if (main_inout_8x4_inout_8x4_override_en) begin
		main_inout_8x4_inout_8x4_oe <= main_inout_8x4_inout_8x4_override_oe;
	end else begin
		main_inout_8x4_inout_8x4_oe <= main_inout_8x4_inout_8x4_oe_k;
	end
	main_inout_8x4_inout_8x4_i_d <= main_inout_8x4_serdes_i0[7];
	main_inout_8x4_inout_8x4_iinterface4_stb <= ((main_inout_8x4_inout_8x4_sample | (main_inout_8x4_inout_8x4_sensitivity[0] & (main_inout_8x4_serdes_i0[7] & (~main_inout_8x4_inout_8x4_i_d)))) | (main_inout_8x4_inout_8x4_sensitivity[1] & ((~main_inout_8x4_serdes_i0[7]) & main_inout_8x4_inout_8x4_i_d)));
	main_inout_8x4_inout_8x4_iinterface4_data <= main_inout_8x4_serdes_i0[7];
	main_inout_8x4_inout_8x4_iinterface4_fine_ts <= main_inout_8x4_inout_8x4_o;
	if ((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0))) begin
		main_inout_8x4_inout_8x4_previous_data <= main_inout_8x4_inout_8x4_ointerface4_data[0];
	end
	if (main_inout_8x4_inout_8x4_override_en) begin
		main_inout_8x4_serdes_o0 <= {8{main_inout_8x4_inout_8x4_override_o}};
	end else begin
		if ((((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0)) & (~main_inout_8x4_inout_8x4_previous_data)) & main_inout_8x4_inout_8x4_ointerface4_data[0])) begin
			main_inout_8x4_serdes_o0 <= builder_sync_f_t_array_muxed16;
		end else begin
			if ((((main_inout_8x4_inout_8x4_ointerface4_stb & (main_inout_8x4_inout_8x4_ointerface4_address == 1'd0)) & main_inout_8x4_inout_8x4_previous_data) & (~main_inout_8x4_inout_8x4_ointerface4_data[0]))) begin
				main_inout_8x4_serdes_o0 <= builder_sync_f_f_array_muxed16;
			end else begin
				main_inout_8x4_serdes_o0 <= {8{main_inout_8x4_inout_8x4_previous_data}};
			end
		end
	end
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd1))) begin
		main_inout_8x5_inout_8x5_oe_k <= main_inout_8x5_inout_8x5_ointerface5_data[0];
	end
	if (main_inout_8x5_inout_8x5_override_en) begin
		main_inout_8x5_inout_8x5_oe <= main_inout_8x5_inout_8x5_override_oe;
	end else begin
		main_inout_8x5_inout_8x5_oe <= main_inout_8x5_inout_8x5_oe_k;
	end
	main_inout_8x5_inout_8x5_i_d <= main_inout_8x5_serdes_i0[7];
	main_inout_8x5_inout_8x5_iinterface5_stb <= ((main_inout_8x5_inout_8x5_sample | (main_inout_8x5_inout_8x5_sensitivity[0] & (main_inout_8x5_serdes_i0[7] & (~main_inout_8x5_inout_8x5_i_d)))) | (main_inout_8x5_inout_8x5_sensitivity[1] & ((~main_inout_8x5_serdes_i0[7]) & main_inout_8x5_inout_8x5_i_d)));
	main_inout_8x5_inout_8x5_iinterface5_data <= main_inout_8x5_serdes_i0[7];
	main_inout_8x5_inout_8x5_iinterface5_fine_ts <= main_inout_8x5_inout_8x5_o;
	if ((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0))) begin
		main_inout_8x5_inout_8x5_previous_data <= main_inout_8x5_inout_8x5_ointerface5_data[0];
	end
	if (main_inout_8x5_inout_8x5_override_en) begin
		main_inout_8x5_serdes_o0 <= {8{main_inout_8x5_inout_8x5_override_o}};
	end else begin
		if ((((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0)) & (~main_inout_8x5_inout_8x5_previous_data)) & main_inout_8x5_inout_8x5_ointerface5_data[0])) begin
			main_inout_8x5_serdes_o0 <= builder_sync_f_t_array_muxed17;
		end else begin
			if ((((main_inout_8x5_inout_8x5_ointerface5_stb & (main_inout_8x5_inout_8x5_ointerface5_address == 1'd0)) & main_inout_8x5_inout_8x5_previous_data) & (~main_inout_8x5_inout_8x5_ointerface5_data[0]))) begin
				main_inout_8x5_serdes_o0 <= builder_sync_f_f_array_muxed17;
			end else begin
				main_inout_8x5_serdes_o0 <= {8{main_inout_8x5_inout_8x5_previous_data}};
			end
		end
	end
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd1))) begin
		main_inout_8x6_inout_8x6_oe_k <= main_inout_8x6_inout_8x6_ointerface6_data[0];
	end
	if (main_inout_8x6_inout_8x6_override_en) begin
		main_inout_8x6_inout_8x6_oe <= main_inout_8x6_inout_8x6_override_oe;
	end else begin
		main_inout_8x6_inout_8x6_oe <= main_inout_8x6_inout_8x6_oe_k;
	end
	main_inout_8x6_inout_8x6_i_d <= main_inout_8x6_serdes_i0[7];
	main_inout_8x6_inout_8x6_iinterface6_stb <= ((main_inout_8x6_inout_8x6_sample | (main_inout_8x6_inout_8x6_sensitivity[0] & (main_inout_8x6_serdes_i0[7] & (~main_inout_8x6_inout_8x6_i_d)))) | (main_inout_8x6_inout_8x6_sensitivity[1] & ((~main_inout_8x6_serdes_i0[7]) & main_inout_8x6_inout_8x6_i_d)));
	main_inout_8x6_inout_8x6_iinterface6_data <= main_inout_8x6_serdes_i0[7];
	main_inout_8x6_inout_8x6_iinterface6_fine_ts <= main_inout_8x6_inout_8x6_o;
	if ((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0))) begin
		main_inout_8x6_inout_8x6_previous_data <= main_inout_8x6_inout_8x6_ointerface6_data[0];
	end
	if (main_inout_8x6_inout_8x6_override_en) begin
		main_inout_8x6_serdes_o0 <= {8{main_inout_8x6_inout_8x6_override_o}};
	end else begin
		if ((((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0)) & (~main_inout_8x6_inout_8x6_previous_data)) & main_inout_8x6_inout_8x6_ointerface6_data[0])) begin
			main_inout_8x6_serdes_o0 <= builder_sync_f_t_array_muxed18;
		end else begin
			if ((((main_inout_8x6_inout_8x6_ointerface6_stb & (main_inout_8x6_inout_8x6_ointerface6_address == 1'd0)) & main_inout_8x6_inout_8x6_previous_data) & (~main_inout_8x6_inout_8x6_ointerface6_data[0]))) begin
				main_inout_8x6_serdes_o0 <= builder_sync_f_f_array_muxed18;
			end else begin
				main_inout_8x6_serdes_o0 <= {8{main_inout_8x6_inout_8x6_previous_data}};
			end
		end
	end
	if (main_output0_stb) begin
		main_output0_pad_k <= main_output0_data;
	end
	if (main_output0_override_en) begin
		main_output0_pad_o <= main_output0_override_o;
	end else begin
		main_output0_pad_o <= main_output0_pad_k;
	end
	if (main_output1_stb) begin
		main_output1_pad_k <= main_output1_data;
	end
	if (main_output1_override_en) begin
		main_output1_pad_o <= main_output1_override_o;
	end else begin
		main_output1_pad_o <= main_output1_pad_k;
	end
	main_clockgen_acc <= (main_clockgen_acc + main_clockgen_ftw);
	if (main_clockgen_stb) begin
		if ((main_clockgen_data != 1'd0)) begin
			main_clockgen_acc <= 24'd8388608;
		end else begin
			main_clockgen_acc <= 1'd0;
		end
	end
	la32_p <= main_clockgen_acc[23];
	if (main_spimaster0_iinterface0_stb) begin
		main_spimaster0_read <= 1'd0;
	end
	if ((main_spimaster0_ointerface0_stb & main_spimaster0_spimachine0_writable)) begin
		if (main_spimaster0_ointerface0_address) begin
			{main_spimaster0_config_cs, main_spimaster0_config_div, main_spimaster0_config_padding, main_spimaster0_config_length, main_spimaster0_config_half_duplex, main_spimaster0_config_lsb_first, main_spimaster0_config_clk_phase, main_spimaster0_config_clk_polarity, main_spimaster0_config_cs_polarity, main_spimaster0_config_input, main_spimaster0_config_end, main_spimaster0_config_offline} <= main_spimaster0_ointerface0_data;
		end else begin
			main_spimaster0_read <= main_spimaster0_config_input;
		end
	end
	if (main_spimaster0_interface_ce) begin
		main_spimaster0_interface_cs_o <= (({1{main_spimaster0_interface_cs_next}} & main_spimaster0_interface_cs) ^ (~main_spimaster0_interface_cs_polarity));
		main_spimaster0_interface_clk_o <= (main_spimaster0_interface_clk_next ^ main_spimaster0_interface_clk_polarity);
	end
	if (main_spimaster0_interface_sample) begin
		main_spimaster0_interface_miso_reg <= main_spimaster0_interface_miso_i;
		main_spimaster0_interface_mosi_reg <= main_spimaster0_interface_mosi_i;
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_n <= main_spimaster0_spimachine0_length;
		main_spimaster0_spimachine0_end1 <= main_spimaster0_spimachine0_end0;
	end
	if (main_spimaster0_spimachine0_shift) begin
		main_spimaster0_spimachine0_n <= (main_spimaster0_spimachine0_n - 1'd1);
	end
	if (main_spimaster0_spimachine0_shift) begin
		main_spimaster0_spimachine0_sr <= main_spimaster0_spimachine0_pdi;
		main_spimaster0_spimachine0_sdo <= (main_spimaster0_spimachine0_lsb_first ? main_spimaster0_spimachine0_pdi[0] : main_spimaster0_spimachine0_pdi[31]);
	end
	if (main_spimaster0_spimachine0_load1) begin
		main_spimaster0_spimachine0_sr <= main_spimaster0_spimachine0_pdo;
		main_spimaster0_spimachine0_sdo <= (main_spimaster0_spimachine0_lsb_first ? main_spimaster0_spimachine0_pdo[0] : main_spimaster0_spimachine0_pdo[31]);
	end
	if (main_spimaster0_spimachine0_count) begin
		if (main_spimaster0_spimachine0_cnt_done) begin
			if (main_spimaster0_spimachine0_do_extend) begin
				main_spimaster0_spimachine0_do_extend <= 1'd0;
			end else begin
				main_spimaster0_spimachine0_cnt <= main_spimaster0_spimachine0_div[7:1];
				main_spimaster0_spimachine0_do_extend <= (main_spimaster0_spimachine0_extend & main_spimaster0_spimachine0_div[0]);
			end
		end else begin
			main_spimaster0_spimachine0_cnt <= (main_spimaster0_spimachine0_cnt - 1'd1);
		end
	end
	builder_spimaster0_state <= builder_spimaster0_next_state;
	if (main_spimaster1_iinterface1_stb) begin
		main_spimaster1_read <= 1'd0;
	end
	if ((main_spimaster1_ointerface1_stb & main_spimaster1_spimachine1_writable)) begin
		if (main_spimaster1_ointerface1_address) begin
			{main_spimaster1_config_cs, main_spimaster1_config_div, main_spimaster1_config_padding, main_spimaster1_config_length, main_spimaster1_config_half_duplex, main_spimaster1_config_lsb_first, main_spimaster1_config_clk_phase, main_spimaster1_config_clk_polarity, main_spimaster1_config_cs_polarity, main_spimaster1_config_input, main_spimaster1_config_end, main_spimaster1_config_offline} <= main_spimaster1_ointerface1_data;
		end else begin
			main_spimaster1_read <= main_spimaster1_config_input;
		end
	end
	if (main_spimaster1_interface_ce) begin
		main_spimaster1_interface_cs_o <= (({1{main_spimaster1_interface_cs_next}} & main_spimaster1_interface_cs) ^ (~main_spimaster1_interface_cs_polarity));
		main_spimaster1_interface_clk_o <= (main_spimaster1_interface_clk_next ^ main_spimaster1_interface_clk_polarity);
	end
	if (main_spimaster1_interface_sample) begin
		main_spimaster1_interface_miso_reg <= main_spimaster1_interface_miso_i;
		main_spimaster1_interface_mosi_reg <= main_spimaster1_interface_mosi_i;
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_n <= main_spimaster1_spimachine1_length;
		main_spimaster1_spimachine1_end1 <= main_spimaster1_spimachine1_end0;
	end
	if (main_spimaster1_spimachine1_shift) begin
		main_spimaster1_spimachine1_n <= (main_spimaster1_spimachine1_n - 1'd1);
	end
	if (main_spimaster1_spimachine1_shift) begin
		main_spimaster1_spimachine1_sr <= main_spimaster1_spimachine1_pdi;
		main_spimaster1_spimachine1_sdo <= (main_spimaster1_spimachine1_lsb_first ? main_spimaster1_spimachine1_pdi[0] : main_spimaster1_spimachine1_pdi[31]);
	end
	if (main_spimaster1_spimachine1_load1) begin
		main_spimaster1_spimachine1_sr <= main_spimaster1_spimachine1_pdo;
		main_spimaster1_spimachine1_sdo <= (main_spimaster1_spimachine1_lsb_first ? main_spimaster1_spimachine1_pdo[0] : main_spimaster1_spimachine1_pdo[31]);
	end
	if (main_spimaster1_spimachine1_count) begin
		if (main_spimaster1_spimachine1_cnt_done) begin
			if (main_spimaster1_spimachine1_do_extend) begin
				main_spimaster1_spimachine1_do_extend <= 1'd0;
			end else begin
				main_spimaster1_spimachine1_cnt <= main_spimaster1_spimachine1_div[7:1];
				main_spimaster1_spimachine1_do_extend <= (main_spimaster1_spimachine1_extend & main_spimaster1_spimachine1_div[0]);
			end
		end else begin
			main_spimaster1_spimachine1_cnt <= (main_spimaster1_spimachine1_cnt - 1'd1);
		end
	end
	builder_spimaster1_state <= builder_spimaster1_next_state;
	if (main_spimaster2_iinterface2_stb) begin
		main_spimaster2_read <= 1'd0;
	end
	if ((main_spimaster2_ointerface2_stb & main_spimaster2_spimachine2_writable)) begin
		if (main_spimaster2_ointerface2_address) begin
			{main_spimaster2_config_cs, main_spimaster2_config_div, main_spimaster2_config_padding, main_spimaster2_config_length, main_spimaster2_config_half_duplex, main_spimaster2_config_lsb_first, main_spimaster2_config_clk_phase, main_spimaster2_config_clk_polarity, main_spimaster2_config_cs_polarity, main_spimaster2_config_input, main_spimaster2_config_end, main_spimaster2_config_offline} <= main_spimaster2_ointerface2_data;
		end else begin
			main_spimaster2_read <= main_spimaster2_config_input;
		end
	end
	if (main_spimaster2_interface_ce) begin
		main_spimaster2_interface_cs_o <= (({1{main_spimaster2_interface_cs_next}} & main_spimaster2_interface_cs) ^ (~main_spimaster2_interface_cs_polarity));
		main_spimaster2_interface_clk_o <= (main_spimaster2_interface_clk_next ^ main_spimaster2_interface_clk_polarity);
	end
	if (main_spimaster2_interface_sample) begin
		main_spimaster2_interface_miso_reg <= main_spimaster2_interface_miso_i;
		main_spimaster2_interface_mosi_reg <= main_spimaster2_interface_mosi_i;
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_n <= main_spimaster2_spimachine2_length;
		main_spimaster2_spimachine2_end1 <= main_spimaster2_spimachine2_end0;
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_n <= (main_spimaster2_spimachine2_n - 1'd1);
	end
	if (main_spimaster2_spimachine2_shift) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdi;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdi[0] : main_spimaster2_spimachine2_pdi[31]);
	end
	if (main_spimaster2_spimachine2_load1) begin
		main_spimaster2_spimachine2_sr <= main_spimaster2_spimachine2_pdo;
		main_spimaster2_spimachine2_sdo <= (main_spimaster2_spimachine2_lsb_first ? main_spimaster2_spimachine2_pdo[0] : main_spimaster2_spimachine2_pdo[31]);
	end
	if (main_spimaster2_spimachine2_count) begin
		if (main_spimaster2_spimachine2_cnt_done) begin
			if (main_spimaster2_spimachine2_do_extend) begin
				main_spimaster2_spimachine2_do_extend <= 1'd0;
			end else begin
				main_spimaster2_spimachine2_cnt <= main_spimaster2_spimachine2_div[7:1];
				main_spimaster2_spimachine2_do_extend <= (main_spimaster2_spimachine2_extend & main_spimaster2_spimachine2_div[0]);
			end
		end else begin
			main_spimaster2_spimachine2_cnt <= (main_spimaster2_spimachine2_cnt - 1'd1);
		end
	end
	builder_spimaster2_state <= builder_spimaster2_next_state;
	if (main_spimaster3_iinterface3_stb) begin
		main_spimaster3_read <= 1'd0;
	end
	if ((main_spimaster3_ointerface3_stb & main_spimaster3_spimachine3_writable)) begin
		if (main_spimaster3_ointerface3_address) begin
			{main_spimaster3_config_cs, main_spimaster3_config_div, main_spimaster3_config_padding, main_spimaster3_config_length, main_spimaster3_config_half_duplex, main_spimaster3_config_lsb_first, main_spimaster3_config_clk_phase, main_spimaster3_config_clk_polarity, main_spimaster3_config_cs_polarity, main_spimaster3_config_input, main_spimaster3_config_end, main_spimaster3_config_offline} <= main_spimaster3_ointerface3_data;
		end else begin
			main_spimaster3_read <= main_spimaster3_config_input;
		end
	end
	if (main_spimaster3_interface_ce) begin
		main_spimaster3_interface_cs_o <= (({1{main_spimaster3_interface_cs_next}} & main_spimaster3_interface_cs) ^ (~main_spimaster3_interface_cs_polarity));
		main_spimaster3_interface_clk_o <= (main_spimaster3_interface_clk_next ^ main_spimaster3_interface_clk_polarity);
	end
	if (main_spimaster3_interface_sample) begin
		main_spimaster3_interface_miso_reg <= main_spimaster3_interface_miso_i;
		main_spimaster3_interface_mosi_reg <= main_spimaster3_interface_mosi_i;
	end
	if (main_spimaster3_spimachine3_load1) begin
		main_spimaster3_spimachine3_n <= main_spimaster3_spimachine3_length;
		main_spimaster3_spimachine3_end1 <= main_spimaster3_spimachine3_end0;
	end
	if (main_spimaster3_spimachine3_shift) begin
		main_spimaster3_spimachine3_n <= (main_spimaster3_spimachine3_n - 1'd1);
	end
	if (main_spimaster3_spimachine3_shift) begin
		main_spimaster3_spimachine3_sr <= main_spimaster3_spimachine3_pdi;
		main_spimaster3_spimachine3_sdo <= (main_spimaster3_spimachine3_lsb_first ? main_spimaster3_spimachine3_pdi[0] : main_spimaster3_spimachine3_pdi[31]);
	end
	if (main_spimaster3_spimachine3_load1) begin
		main_spimaster3_spimachine3_sr <= main_spimaster3_spimachine3_pdo;
		main_spimaster3_spimachine3_sdo <= (main_spimaster3_spimachine3_lsb_first ? main_spimaster3_spimachine3_pdo[0] : main_spimaster3_spimachine3_pdo[31]);
	end
	if (main_spimaster3_spimachine3_count) begin
		if (main_spimaster3_spimachine3_cnt_done) begin
			if (main_spimaster3_spimachine3_do_extend) begin
				main_spimaster3_spimachine3_do_extend <= 1'd0;
			end else begin
				main_spimaster3_spimachine3_cnt <= main_spimaster3_spimachine3_div[7:1];
				main_spimaster3_spimachine3_do_extend <= (main_spimaster3_spimachine3_extend & main_spimaster3_spimachine3_div[0]);
			end
		end else begin
			main_spimaster3_spimachine3_cnt <= (main_spimaster3_spimachine3_cnt - 1'd1);
		end
	end
	builder_spimaster3_state <= builder_spimaster3_next_state;
	if (main_spimaster4_iinterface4_stb) begin
		main_spimaster4_read <= 1'd0;
	end
	if ((main_spimaster4_ointerface4_stb & main_spimaster4_spimachine4_writable)) begin
		if (main_spimaster4_ointerface4_address) begin
			{main_spimaster4_config_cs, main_spimaster4_config_div, main_spimaster4_config_padding, main_spimaster4_config_length, main_spimaster4_config_half_duplex, main_spimaster4_config_lsb_first, main_spimaster4_config_clk_phase, main_spimaster4_config_clk_polarity, main_spimaster4_config_cs_polarity, main_spimaster4_config_input, main_spimaster4_config_end, main_spimaster4_config_offline} <= main_spimaster4_ointerface4_data;
		end else begin
			main_spimaster4_read <= main_spimaster4_config_input;
		end
	end
	if (main_spimaster4_interface_ce) begin
		main_spimaster4_interface_cs_o <= (({1{main_spimaster4_interface_cs_next}} & main_spimaster4_interface_cs) ^ (~main_spimaster4_interface_cs_polarity));
		main_spimaster4_interface_clk_o <= (main_spimaster4_interface_clk_next ^ main_spimaster4_interface_clk_polarity);
	end
	if (main_spimaster4_interface_sample) begin
		main_spimaster4_interface_miso_reg <= main_spimaster4_interface_miso_i;
		main_spimaster4_interface_mosi_reg <= main_spimaster4_interface_mosi_i;
	end
	if (main_spimaster4_spimachine4_load1) begin
		main_spimaster4_spimachine4_n <= main_spimaster4_spimachine4_length;
		main_spimaster4_spimachine4_end1 <= main_spimaster4_spimachine4_end0;
	end
	if (main_spimaster4_spimachine4_shift) begin
		main_spimaster4_spimachine4_n <= (main_spimaster4_spimachine4_n - 1'd1);
	end
	if (main_spimaster4_spimachine4_shift) begin
		main_spimaster4_spimachine4_sr <= main_spimaster4_spimachine4_pdi;
		main_spimaster4_spimachine4_sdo <= (main_spimaster4_spimachine4_lsb_first ? main_spimaster4_spimachine4_pdi[0] : main_spimaster4_spimachine4_pdi[31]);
	end
	if (main_spimaster4_spimachine4_load1) begin
		main_spimaster4_spimachine4_sr <= main_spimaster4_spimachine4_pdo;
		main_spimaster4_spimachine4_sdo <= (main_spimaster4_spimachine4_lsb_first ? main_spimaster4_spimachine4_pdo[0] : main_spimaster4_spimachine4_pdo[31]);
	end
	if (main_spimaster4_spimachine4_count) begin
		if (main_spimaster4_spimachine4_cnt_done) begin
			if (main_spimaster4_spimachine4_do_extend) begin
				main_spimaster4_spimachine4_do_extend <= 1'd0;
			end else begin
				main_spimaster4_spimachine4_cnt <= main_spimaster4_spimachine4_div[7:1];
				main_spimaster4_spimachine4_do_extend <= (main_spimaster4_spimachine4_extend & main_spimaster4_spimachine4_div[0]);
			end
		end else begin
			main_spimaster4_spimachine4_cnt <= (main_spimaster4_spimachine4_cnt - 1'd1);
		end
	end
	builder_spimaster4_state <= builder_spimaster4_next_state;
	if (main_ad9914_current_sel[0]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws0[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws0[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[1]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws1[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws1[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[2]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws2[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws2[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[3]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws3[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws3[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[4]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws4[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws4[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[5]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws5[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws5[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[6]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws6[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws6[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[7]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws7[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws7[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[8]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws8[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws8[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[9]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws9[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws9[31:16] <= main_ad9914_current_data;
		end
	end
	if (main_ad9914_current_sel[10]) begin
		if ((main_ad9914_current_address == 5'd17)) begin
			main_ad9914_ftws10[15:0] <= main_ad9914_current_data;
		end
		if ((main_ad9914_current_address == 5'd19)) begin
			main_ad9914_ftws10[31:16] <= main_ad9914_current_data;
		end
	end
	if ((main_ad9914_current_address == 8'd128)) begin
		if (main_ad9914_current_sel[0]) begin
			main_ad9914_probes0 <= main_ad9914_ftws0;
		end
		if (main_ad9914_current_sel[1]) begin
			main_ad9914_probes1 <= main_ad9914_ftws1;
		end
		if (main_ad9914_current_sel[2]) begin
			main_ad9914_probes2 <= main_ad9914_ftws2;
		end
		if (main_ad9914_current_sel[3]) begin
			main_ad9914_probes3 <= main_ad9914_ftws3;
		end
		if (main_ad9914_current_sel[4]) begin
			main_ad9914_probes4 <= main_ad9914_ftws4;
		end
		if (main_ad9914_current_sel[5]) begin
			main_ad9914_probes5 <= main_ad9914_ftws5;
		end
		if (main_ad9914_current_sel[6]) begin
			main_ad9914_probes6 <= main_ad9914_ftws6;
		end
		if (main_ad9914_current_sel[7]) begin
			main_ad9914_probes7 <= main_ad9914_ftws7;
		end
		if (main_ad9914_current_sel[8]) begin
			main_ad9914_probes8 <= main_ad9914_ftws8;
		end
		if (main_ad9914_current_sel[9]) begin
			main_ad9914_probes9 <= main_ad9914_ftws9;
		end
		if (main_ad9914_current_sel[10]) begin
			main_ad9914_probes10 <= main_ad9914_ftws10;
		end
	end
	if ((~main_ad9914_hold_address)) begin
		dds_a <= main_ad9914_bus_adr;
	end
	main_ad9914_o <= main_ad9914_bus_dat_w;
	main_ad9914_dr <= main_ad9914_i;
	main_ad9914_oe <= (~main_ad9914_rx);
	if (main_ad9914_gpio_load) begin
		main_ad9914_gpio <= main_ad9914_bus_dat_w;
	end
	dds_fud <= main_ad9914_fud;
	dds_wr_n <= (~main_ad9914_wr);
	dds_rd_n <= (~main_ad9914_rd);
	if (main_ad9914_read_timer_wait) begin
		if ((~main_ad9914_read_timer_done)) begin
			main_ad9914_read_timer_count <= (main_ad9914_read_timer_count - 1'd1);
		end
	end else begin
		main_ad9914_read_timer_count <= 4'd10;
	end
	if (main_ad9914_hiz_timer_wait) begin
		if ((~main_ad9914_hiz_timer_done)) begin
			main_ad9914_hiz_timer_count <= (main_ad9914_hiz_timer_count - 1'd1);
		end
	end else begin
		main_ad9914_hiz_timer_count <= 2'd3;
	end
	builder_ad9914_state <= builder_ad9914_next_state;
	if (rio_phy_rst) begin
		main_output_8x0_o <= 8'd0;
		main_output_8x0_previous_data <= 1'd0;
		main_output_8x1_o <= 8'd0;
		main_output_8x1_previous_data <= 1'd0;
		main_output_8x2_o <= 8'd0;
		main_output_8x2_previous_data <= 1'd0;
		main_inout_8x0_serdes_o0 <= 8'd0;
		main_inout_8x0_inout_8x0_iinterface0_stb <= 1'd0;
		main_inout_8x0_inout_8x0_oe <= 1'd0;
		main_inout_8x0_inout_8x0_previous_data <= 1'd0;
		main_inout_8x0_inout_8x0_oe_k <= 1'd0;
		main_inout_8x0_inout_8x0_i_d <= 1'd0;
		main_output_8x3_o <= 8'd0;
		main_output_8x3_previous_data <= 1'd0;
		main_output_8x4_o <= 8'd0;
		main_output_8x4_previous_data <= 1'd0;
		main_output_8x5_o <= 8'd0;
		main_output_8x5_previous_data <= 1'd0;
		main_inout_8x1_serdes_o0 <= 8'd0;
		main_inout_8x1_inout_8x1_iinterface1_stb <= 1'd0;
		main_inout_8x1_inout_8x1_oe <= 1'd0;
		main_inout_8x1_inout_8x1_previous_data <= 1'd0;
		main_inout_8x1_inout_8x1_oe_k <= 1'd0;
		main_inout_8x1_inout_8x1_i_d <= 1'd0;
		main_output_8x6_o <= 8'd0;
		main_output_8x6_previous_data <= 1'd0;
		main_output_8x7_o <= 8'd0;
		main_output_8x7_previous_data <= 1'd0;
		main_output_8x8_o <= 8'd0;
		main_output_8x8_previous_data <= 1'd0;
		main_inout_8x2_serdes_o0 <= 8'd0;
		main_inout_8x2_inout_8x2_iinterface2_stb <= 1'd0;
		main_inout_8x2_inout_8x2_oe <= 1'd0;
		main_inout_8x2_inout_8x2_previous_data <= 1'd0;
		main_inout_8x2_inout_8x2_oe_k <= 1'd0;
		main_inout_8x2_inout_8x2_i_d <= 1'd0;
		main_output_8x9_o <= 8'd0;
		main_output_8x9_previous_data <= 1'd0;
		main_output_8x10_o <= 8'd0;
		main_output_8x10_previous_data <= 1'd0;
		main_output_8x11_o <= 8'd0;
		main_output_8x11_previous_data <= 1'd0;
		main_inout_8x3_serdes_o0 <= 8'd0;
		main_inout_8x3_inout_8x3_iinterface3_stb <= 1'd0;
		main_inout_8x3_inout_8x3_oe <= 1'd0;
		main_inout_8x3_inout_8x3_previous_data <= 1'd0;
		main_inout_8x3_inout_8x3_oe_k <= 1'd0;
		main_inout_8x3_inout_8x3_i_d <= 1'd0;
		main_inout_8x4_serdes_o0 <= 8'd0;
		main_inout_8x4_inout_8x4_iinterface4_stb <= 1'd0;
		main_inout_8x4_inout_8x4_oe <= 1'd0;
		main_inout_8x4_inout_8x4_previous_data <= 1'd0;
		main_inout_8x4_inout_8x4_oe_k <= 1'd0;
		main_inout_8x4_inout_8x4_i_d <= 1'd0;
		main_inout_8x5_serdes_o0 <= 8'd0;
		main_inout_8x5_inout_8x5_iinterface5_stb <= 1'd0;
		main_inout_8x5_inout_8x5_oe <= 1'd0;
		main_inout_8x5_inout_8x5_previous_data <= 1'd0;
		main_inout_8x5_inout_8x5_oe_k <= 1'd0;
		main_inout_8x5_inout_8x5_i_d <= 1'd0;
		main_inout_8x6_serdes_o0 <= 8'd0;
		main_inout_8x6_inout_8x6_iinterface6_stb <= 1'd0;
		main_inout_8x6_inout_8x6_oe <= 1'd0;
		main_inout_8x6_inout_8x6_previous_data <= 1'd0;
		main_inout_8x6_inout_8x6_oe_k <= 1'd0;
		main_inout_8x6_inout_8x6_i_d <= 1'd0;
		main_output0_pad_k <= 1'd0;
		main_output1_pad_k <= 1'd0;
		la32_p <= 1'd0;
		main_clockgen_acc <= 24'd0;
		main_spimaster0_interface_cs_o <= 1'd1;
		main_spimaster0_interface_clk_o <= 1'd0;
		main_spimaster0_spimachine0_cnt <= 7'd0;
		main_spimaster0_spimachine0_do_extend <= 1'd0;
		main_spimaster0_config_offline <= 1'd1;
		main_spimaster0_config_end <= 1'd1;
		main_spimaster0_config_input <= 1'd0;
		main_spimaster0_config_cs_polarity <= 1'd0;
		main_spimaster0_config_clk_polarity <= 1'd0;
		main_spimaster0_config_clk_phase <= 1'd0;
		main_spimaster0_config_lsb_first <= 1'd0;
		main_spimaster0_config_half_duplex <= 1'd0;
		main_spimaster0_config_length <= 5'd0;
		main_spimaster0_config_padding <= 3'd0;
		main_spimaster0_config_div <= 8'd0;
		main_spimaster0_config_cs <= 8'd0;
		main_spimaster0_read <= 1'd0;
		main_spimaster1_interface_cs_o <= 1'd1;
		main_spimaster1_interface_clk_o <= 1'd0;
		main_spimaster1_spimachine1_cnt <= 7'd0;
		main_spimaster1_spimachine1_do_extend <= 1'd0;
		main_spimaster1_config_offline <= 1'd1;
		main_spimaster1_config_end <= 1'd1;
		main_spimaster1_config_input <= 1'd0;
		main_spimaster1_config_cs_polarity <= 1'd0;
		main_spimaster1_config_clk_polarity <= 1'd0;
		main_spimaster1_config_clk_phase <= 1'd0;
		main_spimaster1_config_lsb_first <= 1'd0;
		main_spimaster1_config_half_duplex <= 1'd0;
		main_spimaster1_config_length <= 5'd0;
		main_spimaster1_config_padding <= 3'd0;
		main_spimaster1_config_div <= 8'd0;
		main_spimaster1_config_cs <= 8'd0;
		main_spimaster1_read <= 1'd0;
		main_spimaster2_interface_cs_o <= 1'd1;
		main_spimaster2_interface_clk_o <= 1'd0;
		main_spimaster2_spimachine2_cnt <= 7'd0;
		main_spimaster2_spimachine2_do_extend <= 1'd0;
		main_spimaster2_config_offline <= 1'd1;
		main_spimaster2_config_end <= 1'd1;
		main_spimaster2_config_input <= 1'd0;
		main_spimaster2_config_cs_polarity <= 1'd0;
		main_spimaster2_config_clk_polarity <= 1'd0;
		main_spimaster2_config_clk_phase <= 1'd0;
		main_spimaster2_config_lsb_first <= 1'd0;
		main_spimaster2_config_half_duplex <= 1'd0;
		main_spimaster2_config_length <= 5'd0;
		main_spimaster2_config_padding <= 3'd0;
		main_spimaster2_config_div <= 8'd0;
		main_spimaster2_config_cs <= 8'd0;
		main_spimaster2_read <= 1'd0;
		main_spimaster3_interface_cs_o <= 1'd1;
		main_spimaster3_interface_clk_o <= 1'd0;
		main_spimaster3_spimachine3_cnt <= 7'd0;
		main_spimaster3_spimachine3_do_extend <= 1'd0;
		main_spimaster3_config_offline <= 1'd1;
		main_spimaster3_config_end <= 1'd1;
		main_spimaster3_config_input <= 1'd0;
		main_spimaster3_config_cs_polarity <= 1'd0;
		main_spimaster3_config_clk_polarity <= 1'd0;
		main_spimaster3_config_clk_phase <= 1'd0;
		main_spimaster3_config_lsb_first <= 1'd0;
		main_spimaster3_config_half_duplex <= 1'd0;
		main_spimaster3_config_length <= 5'd0;
		main_spimaster3_config_padding <= 3'd0;
		main_spimaster3_config_div <= 8'd0;
		main_spimaster3_config_cs <= 8'd0;
		main_spimaster3_read <= 1'd0;
		main_spimaster4_interface_cs_o <= 1'd1;
		main_spimaster4_interface_clk_o <= 1'd0;
		main_spimaster4_spimachine4_cnt <= 7'd0;
		main_spimaster4_spimachine4_do_extend <= 1'd0;
		main_spimaster4_config_offline <= 1'd1;
		main_spimaster4_config_end <= 1'd1;
		main_spimaster4_config_input <= 1'd0;
		main_spimaster4_config_cs_polarity <= 1'd0;
		main_spimaster4_config_clk_polarity <= 1'd0;
		main_spimaster4_config_clk_phase <= 1'd0;
		main_spimaster4_config_lsb_first <= 1'd0;
		main_spimaster4_config_half_duplex <= 1'd0;
		main_spimaster4_config_length <= 5'd0;
		main_spimaster4_config_padding <= 3'd0;
		main_spimaster4_config_div <= 8'd0;
		main_spimaster4_config_cs <= 8'd0;
		main_spimaster4_read <= 1'd0;
		dds_a <= 7'd0;
		dds_fud <= 1'd0;
		dds_wr_n <= 1'd1;
		dds_rd_n <= 1'd1;
		main_ad9914_o <= 16'd0;
		main_ad9914_oe <= 1'd0;
		main_ad9914_dr <= 16'd0;
		main_ad9914_gpio <= 12'd0;
		main_ad9914_read_timer_count <= 4'd10;
		main_ad9914_hiz_timer_count <= 2'd3;
		main_ad9914_probes0 <= 32'd0;
		main_ad9914_probes1 <= 32'd0;
		main_ad9914_probes2 <= 32'd0;
		main_ad9914_probes3 <= 32'd0;
		main_ad9914_probes4 <= 32'd0;
		main_ad9914_probes5 <= 32'd0;
		main_ad9914_probes6 <= 32'd0;
		main_ad9914_probes7 <= 32'd0;
		main_ad9914_probes8 <= 32'd0;
		main_ad9914_probes9 <= 32'd0;
		main_ad9914_probes10 <= 32'd0;
		main_ad9914_ftws0 <= 32'd0;
		main_ad9914_ftws1 <= 32'd0;
		main_ad9914_ftws2 <= 32'd0;
		main_ad9914_ftws3 <= 32'd0;
		main_ad9914_ftws4 <= 32'd0;
		main_ad9914_ftws5 <= 32'd0;
		main_ad9914_ftws6 <= 32'd0;
		main_ad9914_ftws7 <= 32'd0;
		main_ad9914_ftws8 <= 32'd0;
		main_ad9914_ftws9 <= 32'd0;
		main_ad9914_ftws10 <= 32'd0;
		builder_spimaster0_state <= 3'd0;
		builder_spimaster1_state <= 3'd0;
		builder_spimaster2_state <= 3'd0;
		builder_spimaster3_state <= 3'd0;
		builder_spimaster4_state <= 3'd0;
		builder_ad9914_state <= 3'd0;
	end
end

always @(posedge rsys_clk) begin
	main_rtio_core_outputs_lanedistributor_min_minus_timestamp <= (main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_laneAmin_minus_timestamp <= (builder_sync_rhs_array_muxed0 - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_laneBmin_minus_timestamp <= (builder_sync_rhs_array_muxed1 - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_last_minus_timestamp <= (main_rtio_core_outputs_lanedistributor_last_coarse_timestamp - main_rtio_core_outputs_lanedistributor_coarse_timestamp);
	main_rtio_core_outputs_lanedistributor_quash <= 1'd0;
	if ((main_rtio_core_cri_chan_sel[15:0] == 5'd28)) begin
		main_rtio_core_outputs_lanedistributor_quash <= 1'd1;
	end
	if (main_rtio_core_outputs_lanedistributor_do_write) begin
		main_rtio_core_outputs_lanedistributor_current_lane <= main_rtio_core_outputs_lanedistributor_use_lanen;
		main_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= main_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		builder_sync_t_lhs_array_muxed = main_rtio_core_outputs_lanedistributor_compensated_timestamp[63:3];
		case (main_rtio_core_outputs_lanedistributor_use_lanen)
			1'd0: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= builder_sync_t_lhs_array_muxed;
			end
			1'd1: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= builder_sync_t_lhs_array_muxed;
			end
			2'd2: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= builder_sync_t_lhs_array_muxed;
			end
			2'd3: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= builder_sync_t_lhs_array_muxed;
			end
			3'd4: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= builder_sync_t_lhs_array_muxed;
			end
			3'd5: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= builder_sync_t_lhs_array_muxed;
			end
			3'd6: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= builder_sync_t_lhs_array_muxed;
			end
			default: begin
				main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= builder_sync_t_lhs_array_muxed;
			end
		endcase
		main_rtio_core_outputs_lanedistributor_seqn <= (main_rtio_core_outputs_lanedistributor_seqn + 1'd1);
	end
	if ((main_rtio_core_cri_cmd == 1'd1)) begin
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
	end
	if (main_rtio_core_outputs_lanedistributor_do_underflow) begin
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd1;
	end
	main_rtio_core_outputs_lanedistributor_sequence_error <= main_rtio_core_outputs_lanedistributor_do_sequence_error;
	main_rtio_core_outputs_lanedistributor_sequence_error_channel <= main_rtio_core_cri_chan_sel[15:0];
	main_rtio_core_outputs_lanedistributor_current_lane_writable_r <= main_rtio_core_outputs_lanedistributor_current_lane_writable;
	if (((~main_rtio_core_outputs_lanedistributor_current_lane_writable_r) & main_rtio_core_outputs_lanedistributor_current_lane_writable)) begin
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd1;
	end
	if (main_rtio_core_outputs_lanedistributor_do_write) begin
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
	end
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_next;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_next;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_next;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_next;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_next;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_next;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_next;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next_binary;
	main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_next;
	if ((main_rtio_core_inputs_selected0 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow0 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer0_o) begin
		main_rtio_core_inputs_overflow0 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected1 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow1 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer1_o) begin
		main_rtio_core_inputs_overflow1 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected2 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow2 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer2_o) begin
		main_rtio_core_inputs_overflow2 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected3 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow3 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer3_o) begin
		main_rtio_core_inputs_overflow3 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected4 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow4 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer4_o) begin
		main_rtio_core_inputs_overflow4 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected5 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow5 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer5_o) begin
		main_rtio_core_inputs_overflow5 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected6 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow6 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer6_o) begin
		main_rtio_core_inputs_overflow6 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected7 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow7 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer7_o) begin
		main_rtio_core_inputs_overflow7 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected8 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow8 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer8_o) begin
		main_rtio_core_inputs_overflow8 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected9 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow9 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer9_o) begin
		main_rtio_core_inputs_overflow9 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected10 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow10 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer10_o) begin
		main_rtio_core_inputs_overflow10 <= 1'd1;
	end
	if ((main_rtio_core_inputs_selected11 & main_rtio_core_inputs_i_ack)) begin
		main_rtio_core_inputs_overflow11 <= 1'd0;
	end
	if (main_rtio_core_inputs_blindtransfer11_o) begin
		main_rtio_core_inputs_overflow11 <= 1'd1;
	end
	main_rtio_core_inputs_i_ack <= 1'd0;
	if (main_rtio_core_inputs_i_ack) begin
		main_rtio_core_cri_i_status <= {1'd0, main_rtio_core_inputs_i_status_raw[1], (~main_rtio_core_inputs_i_status_raw[0])};
		main_rtio_core_cri_i_data <= builder_sync_t_rhs_array_muxed0;
		main_rtio_core_cri_i_timestamp <= builder_sync_t_rhs_array_muxed1;
	end
	if (((main_full_ts_sys >= main_rtio_core_inputs_input_timeout) | (main_rtio_core_inputs_i_status_raw != 1'd0))) begin
		if (main_rtio_core_inputs_input_pending) begin
			main_rtio_core_inputs_i_ack <= 1'd1;
		end
		main_rtio_core_inputs_input_pending <= 1'd0;
	end
	if ((main_rtio_core_cri_cmd == 2'd2)) begin
		main_rtio_core_inputs_input_timeout <= main_rtio_core_cri_i_timeout;
		main_rtio_core_inputs_input_pending <= 1'd1;
		main_rtio_core_cri_i_status <= 3'd4;
	end
	main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_next_binary;
	main_rtio_core_inputs_asyncfifo0_graycounter1_q <= main_rtio_core_inputs_asyncfifo0_graycounter1_q_next;
	main_rtio_core_inputs_blindtransfer0_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer0_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer0_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer0_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_next_binary;
	main_rtio_core_inputs_asyncfifo1_graycounter3_q <= main_rtio_core_inputs_asyncfifo1_graycounter3_q_next;
	main_rtio_core_inputs_blindtransfer1_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer1_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer1_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer1_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_next_binary;
	main_rtio_core_inputs_asyncfifo2_graycounter5_q <= main_rtio_core_inputs_asyncfifo2_graycounter5_q_next;
	main_rtio_core_inputs_blindtransfer2_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer2_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer2_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer2_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_next_binary;
	main_rtio_core_inputs_asyncfifo3_graycounter7_q <= main_rtio_core_inputs_asyncfifo3_graycounter7_q_next;
	main_rtio_core_inputs_blindtransfer3_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer3_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer3_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer3_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_next_binary;
	main_rtio_core_inputs_asyncfifo4_graycounter9_q <= main_rtio_core_inputs_asyncfifo4_graycounter9_q_next;
	main_rtio_core_inputs_blindtransfer4_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer4_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer4_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer4_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_next_binary;
	main_rtio_core_inputs_asyncfifo5_graycounter11_q <= main_rtio_core_inputs_asyncfifo5_graycounter11_q_next;
	main_rtio_core_inputs_blindtransfer5_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer5_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer5_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer5_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_next_binary;
	main_rtio_core_inputs_asyncfifo6_graycounter13_q <= main_rtio_core_inputs_asyncfifo6_graycounter13_q_next;
	main_rtio_core_inputs_blindtransfer6_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer6_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer6_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer6_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_next_binary;
	main_rtio_core_inputs_asyncfifo7_graycounter15_q <= main_rtio_core_inputs_asyncfifo7_graycounter15_q_next;
	main_rtio_core_inputs_blindtransfer7_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer7_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer7_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer7_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_next_binary;
	main_rtio_core_inputs_asyncfifo8_graycounter17_q <= main_rtio_core_inputs_asyncfifo8_graycounter17_q_next;
	main_rtio_core_inputs_blindtransfer8_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer8_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer8_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer8_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_next_binary;
	main_rtio_core_inputs_asyncfifo9_graycounter19_q <= main_rtio_core_inputs_asyncfifo9_graycounter19_q_next;
	main_rtio_core_inputs_blindtransfer9_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer9_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer9_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer9_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_next_binary;
	main_rtio_core_inputs_asyncfifo10_graycounter21_q <= main_rtio_core_inputs_asyncfifo10_graycounter21_q_next;
	main_rtio_core_inputs_blindtransfer10_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer10_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer10_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer10_ps_ack_toggle_i);
	end
	main_rtio_core_inputs_asyncfifo11_graycounter23_q_binary <= main_rtio_core_inputs_asyncfifo11_graycounter23_q_next_binary;
	main_rtio_core_inputs_asyncfifo11_graycounter23_q <= main_rtio_core_inputs_asyncfifo11_graycounter23_q_next;
	main_rtio_core_inputs_blindtransfer11_ps_toggle_o_r <= main_rtio_core_inputs_blindtransfer11_ps_toggle_o;
	if (main_rtio_core_inputs_blindtransfer11_ps_ack_i) begin
		main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_i <= (~main_rtio_core_inputs_blindtransfer11_ps_ack_toggle_i);
	end
	main_rtio_core_o_collision_sync_ps_toggle_o_r <= main_rtio_core_o_collision_sync_ps_toggle_o;
	if (main_rtio_core_o_collision_sync_ps_ack_i) begin
		main_rtio_core_o_collision_sync_ps_ack_toggle_i <= (~main_rtio_core_o_collision_sync_ps_ack_toggle_i);
	end
	main_rtio_core_o_busy_sync_ps_toggle_o_r <= main_rtio_core_o_busy_sync_ps_toggle_o;
	if (main_rtio_core_o_busy_sync_ps_ack_i) begin
		main_rtio_core_o_busy_sync_ps_ack_toggle_i <= (~main_rtio_core_o_busy_sync_ps_ack_toggle_i);
	end
	if (rsys_rst) begin
		main_rtio_core_cri_i_status <= 4'd0;
		main_rtio_core_outputs_lanedistributor_sequence_error <= 1'd0;
		main_rtio_core_outputs_lanedistributor_o_status_underflow <= 1'd0;
		main_rtio_core_outputs_lanedistributor_current_lane <= 3'd0;
		main_rtio_core_outputs_lanedistributor_last_coarse_timestamp <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps0 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps1 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps2 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps3 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps4 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps5 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps6 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_last_lane_coarse_timestamps7 <= 61'd0;
		main_rtio_core_outputs_lanedistributor_seqn <= 12'd0;
		main_rtio_core_outputs_lanedistributor_quash <= 1'd0;
		main_rtio_core_outputs_lanedistributor_force_laneB <= 1'd0;
		main_rtio_core_outputs_lanedistributor_current_lane_writable_r <= 1'd1;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered0_graycounter0_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered1_graycounter2_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered2_graycounter4_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered3_graycounter6_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered4_graycounter8_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered5_graycounter10_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered6_graycounter12_q_binary <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q <= 8'd0;
		main_rtio_core_outputs_asyncfifobuffered7_graycounter14_q_binary <= 8'd0;
		main_rtio_core_inputs_i_ack <= 1'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter1_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo0_graycounter1_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow0 <= 1'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter3_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo1_graycounter3_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow1 <= 1'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter5_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo2_graycounter5_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow2 <= 1'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter7_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo3_graycounter7_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow3 <= 1'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter9_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo4_graycounter9_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow4 <= 1'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter11_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo5_graycounter11_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow5 <= 1'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter13_q <= 10'd0;
		main_rtio_core_inputs_asyncfifo6_graycounter13_q_binary <= 10'd0;
		main_rtio_core_inputs_overflow6 <= 1'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter15_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo7_graycounter15_q_binary <= 3'd0;
		main_rtio_core_inputs_overflow7 <= 1'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter17_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo8_graycounter17_q_binary <= 8'd0;
		main_rtio_core_inputs_overflow8 <= 1'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter19_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo9_graycounter19_q_binary <= 8'd0;
		main_rtio_core_inputs_overflow9 <= 1'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter21_q <= 8'd0;
		main_rtio_core_inputs_asyncfifo10_graycounter21_q_binary <= 8'd0;
		main_rtio_core_inputs_overflow10 <= 1'd0;
		main_rtio_core_inputs_asyncfifo11_graycounter23_q <= 3'd0;
		main_rtio_core_inputs_asyncfifo11_graycounter23_q_binary <= 3'd0;
		main_rtio_core_inputs_overflow11 <= 1'd0;
		main_rtio_core_inputs_input_pending <= 1'd0;
	end
	builder_xilinxmultiregimpl13_regs0 <= main_rtio_core_outputs_asyncfifobuffered0_graycounter1_q;
	builder_xilinxmultiregimpl13_regs1 <= builder_xilinxmultiregimpl13_regs0;
	builder_xilinxmultiregimpl15_regs0 <= main_rtio_core_outputs_asyncfifobuffered1_graycounter3_q;
	builder_xilinxmultiregimpl15_regs1 <= builder_xilinxmultiregimpl15_regs0;
	builder_xilinxmultiregimpl17_regs0 <= main_rtio_core_outputs_asyncfifobuffered2_graycounter5_q;
	builder_xilinxmultiregimpl17_regs1 <= builder_xilinxmultiregimpl17_regs0;
	builder_xilinxmultiregimpl19_regs0 <= main_rtio_core_outputs_asyncfifobuffered3_graycounter7_q;
	builder_xilinxmultiregimpl19_regs1 <= builder_xilinxmultiregimpl19_regs0;
	builder_xilinxmultiregimpl21_regs0 <= main_rtio_core_outputs_asyncfifobuffered4_graycounter9_q;
	builder_xilinxmultiregimpl21_regs1 <= builder_xilinxmultiregimpl21_regs0;
	builder_xilinxmultiregimpl23_regs0 <= main_rtio_core_outputs_asyncfifobuffered5_graycounter11_q;
	builder_xilinxmultiregimpl23_regs1 <= builder_xilinxmultiregimpl23_regs0;
	builder_xilinxmultiregimpl25_regs0 <= main_rtio_core_outputs_asyncfifobuffered6_graycounter13_q;
	builder_xilinxmultiregimpl25_regs1 <= builder_xilinxmultiregimpl25_regs0;
	builder_xilinxmultiregimpl27_regs0 <= main_rtio_core_outputs_asyncfifobuffered7_graycounter15_q;
	builder_xilinxmultiregimpl27_regs1 <= builder_xilinxmultiregimpl27_regs0;
	builder_xilinxmultiregimpl28_regs0 <= main_rtio_core_inputs_asyncfifo0_graycounter0_q;
	builder_xilinxmultiregimpl28_regs1 <= builder_xilinxmultiregimpl28_regs0;
	builder_xilinxmultiregimpl30_regs0 <= main_rtio_core_inputs_blindtransfer0_ps_toggle_i;
	builder_xilinxmultiregimpl30_regs1 <= builder_xilinxmultiregimpl30_regs0;
	builder_xilinxmultiregimpl32_regs0 <= main_rtio_core_inputs_asyncfifo1_graycounter2_q;
	builder_xilinxmultiregimpl32_regs1 <= builder_xilinxmultiregimpl32_regs0;
	builder_xilinxmultiregimpl34_regs0 <= main_rtio_core_inputs_blindtransfer1_ps_toggle_i;
	builder_xilinxmultiregimpl34_regs1 <= builder_xilinxmultiregimpl34_regs0;
	builder_xilinxmultiregimpl36_regs0 <= main_rtio_core_inputs_asyncfifo2_graycounter4_q;
	builder_xilinxmultiregimpl36_regs1 <= builder_xilinxmultiregimpl36_regs0;
	builder_xilinxmultiregimpl38_regs0 <= main_rtio_core_inputs_blindtransfer2_ps_toggle_i;
	builder_xilinxmultiregimpl38_regs1 <= builder_xilinxmultiregimpl38_regs0;
	builder_xilinxmultiregimpl40_regs0 <= main_rtio_core_inputs_asyncfifo3_graycounter6_q;
	builder_xilinxmultiregimpl40_regs1 <= builder_xilinxmultiregimpl40_regs0;
	builder_xilinxmultiregimpl42_regs0 <= main_rtio_core_inputs_blindtransfer3_ps_toggle_i;
	builder_xilinxmultiregimpl42_regs1 <= builder_xilinxmultiregimpl42_regs0;
	builder_xilinxmultiregimpl44_regs0 <= main_rtio_core_inputs_asyncfifo4_graycounter8_q;
	builder_xilinxmultiregimpl44_regs1 <= builder_xilinxmultiregimpl44_regs0;
	builder_xilinxmultiregimpl46_regs0 <= main_rtio_core_inputs_blindtransfer4_ps_toggle_i;
	builder_xilinxmultiregimpl46_regs1 <= builder_xilinxmultiregimpl46_regs0;
	builder_xilinxmultiregimpl48_regs0 <= main_rtio_core_inputs_asyncfifo5_graycounter10_q;
	builder_xilinxmultiregimpl48_regs1 <= builder_xilinxmultiregimpl48_regs0;
	builder_xilinxmultiregimpl50_regs0 <= main_rtio_core_inputs_blindtransfer5_ps_toggle_i;
	builder_xilinxmultiregimpl50_regs1 <= builder_xilinxmultiregimpl50_regs0;
	builder_xilinxmultiregimpl52_regs0 <= main_rtio_core_inputs_asyncfifo6_graycounter12_q;
	builder_xilinxmultiregimpl52_regs1 <= builder_xilinxmultiregimpl52_regs0;
	builder_xilinxmultiregimpl54_regs0 <= main_rtio_core_inputs_blindtransfer6_ps_toggle_i;
	builder_xilinxmultiregimpl54_regs1 <= builder_xilinxmultiregimpl54_regs0;
	builder_xilinxmultiregimpl56_regs0 <= main_rtio_core_inputs_asyncfifo7_graycounter14_q;
	builder_xilinxmultiregimpl56_regs1 <= builder_xilinxmultiregimpl56_regs0;
	builder_xilinxmultiregimpl58_regs0 <= main_rtio_core_inputs_blindtransfer7_ps_toggle_i;
	builder_xilinxmultiregimpl58_regs1 <= builder_xilinxmultiregimpl58_regs0;
	builder_xilinxmultiregimpl60_regs0 <= main_rtio_core_inputs_asyncfifo8_graycounter16_q;
	builder_xilinxmultiregimpl60_regs1 <= builder_xilinxmultiregimpl60_regs0;
	builder_xilinxmultiregimpl62_regs0 <= main_rtio_core_inputs_blindtransfer8_ps_toggle_i;
	builder_xilinxmultiregimpl62_regs1 <= builder_xilinxmultiregimpl62_regs0;
	builder_xilinxmultiregimpl64_regs0 <= main_rtio_core_inputs_asyncfifo9_graycounter18_q;
	builder_xilinxmultiregimpl64_regs1 <= builder_xilinxmultiregimpl64_regs0;
	builder_xilinxmultiregimpl66_regs0 <= main_rtio_core_inputs_blindtransfer9_ps_toggle_i;
	builder_xilinxmultiregimpl66_regs1 <= builder_xilinxmultiregimpl66_regs0;
	builder_xilinxmultiregimpl68_regs0 <= main_rtio_core_inputs_asyncfifo10_graycounter20_q;
	builder_xilinxmultiregimpl68_regs1 <= builder_xilinxmultiregimpl68_regs0;
	builder_xilinxmultiregimpl70_regs0 <= main_rtio_core_inputs_blindtransfer10_ps_toggle_i;
	builder_xilinxmultiregimpl70_regs1 <= builder_xilinxmultiregimpl70_regs0;
	builder_xilinxmultiregimpl72_regs0 <= main_rtio_core_inputs_asyncfifo11_graycounter22_q;
	builder_xilinxmultiregimpl72_regs1 <= builder_xilinxmultiregimpl72_regs0;
	builder_xilinxmultiregimpl74_regs0 <= main_rtio_core_inputs_blindtransfer11_ps_toggle_i;
	builder_xilinxmultiregimpl74_regs1 <= builder_xilinxmultiregimpl74_regs0;
	builder_xilinxmultiregimpl76_regs0 <= main_rtio_core_o_collision_sync_ps_toggle_i;
	builder_xilinxmultiregimpl76_regs1 <= builder_xilinxmultiregimpl76_regs0;
	builder_xilinxmultiregimpl78_regs0 <= main_rtio_core_o_collision_sync_bxfer_data;
	builder_xilinxmultiregimpl78_regs1 <= builder_xilinxmultiregimpl78_regs0;
	builder_xilinxmultiregimpl79_regs0 <= main_rtio_core_o_busy_sync_ps_toggle_i;
	builder_xilinxmultiregimpl79_regs1 <= builder_xilinxmultiregimpl79_regs0;
	builder_xilinxmultiregimpl81_regs0 <= main_rtio_core_o_busy_sync_bxfer_data;
	builder_xilinxmultiregimpl81_regs1 <= builder_xilinxmultiregimpl81_regs0;
end

always @(posedge rtio_clk) begin
	if (main_load) begin
		main_coarse_ts <= main_load_value;
	end else begin
		main_coarse_ts <= (main_coarse_ts + 1'd1);
	end
	main_value_gray_rtio <= (main_i ^ main_i[60:1]);
	if (rtio_rst) begin
		main_coarse_ts <= 61'd0;
	end
end

always @(posedge sys_clk) begin
	main_nist_clock_nist_clock_tmpu_error <= 1'd0;
	if ((main_nist_clock_nist_clock_tmpu_enable_null_storage & (main_nist_clock_nist_clock_dbus_adr[29:10] == 1'd0))) begin
		main_nist_clock_nist_clock_tmpu_error <= 1'd1;
	end
	if ((main_nist_clock_nist_clock_tmpu_enable_prog_storage & (main_nist_clock_nist_clock_dbus_adr[29:10] == main_nist_clock_nist_clock_tmpu_prog_address_storage))) begin
		main_nist_clock_nist_clock_tmpu_error <= 1'd1;
	end
	main_nist_clock_nist_clock_sram_bus_ack <= 1'd0;
	if (((main_nist_clock_nist_clock_sram_bus_cyc & main_nist_clock_nist_clock_sram_bus_stb) & (~main_nist_clock_nist_clock_sram_bus_ack))) begin
		main_nist_clock_nist_clock_sram_bus_ack <= 1'd1;
	end
	main_nist_clock_nist_clock_interface_we <= 1'd0;
	main_nist_clock_nist_clock_interface_dat_w <= main_nist_clock_nist_clock_bus_wishbone_dat_w;
	main_nist_clock_nist_clock_interface_adr <= main_nist_clock_nist_clock_bus_wishbone_adr;
	main_nist_clock_nist_clock_bus_wishbone_dat_r <= main_nist_clock_nist_clock_interface_dat_r;
	if ((main_nist_clock_nist_clock_counter == 1'd1)) begin
		main_nist_clock_nist_clock_interface_we <= main_nist_clock_nist_clock_bus_wishbone_we;
	end
	if ((main_nist_clock_nist_clock_counter == 2'd2)) begin
		main_nist_clock_nist_clock_bus_wishbone_ack <= 1'd1;
	end
	if ((main_nist_clock_nist_clock_counter == 2'd3)) begin
		main_nist_clock_nist_clock_bus_wishbone_ack <= 1'd0;
	end
	if ((main_nist_clock_nist_clock_counter != 1'd0)) begin
		main_nist_clock_nist_clock_counter <= (main_nist_clock_nist_clock_counter + 1'd1);
	end else begin
		if ((main_nist_clock_nist_clock_bus_wishbone_cyc & main_nist_clock_nist_clock_bus_wishbone_stb)) begin
			main_nist_clock_nist_clock_counter <= 1'd1;
		end
	end
	main_nist_clock_nist_clock_uart_phy_sink_ack <= 1'd0;
	if (((main_nist_clock_nist_clock_uart_phy_sink_stb & (~main_nist_clock_nist_clock_uart_phy_tx_busy)) & (~main_nist_clock_nist_clock_uart_phy_sink_ack))) begin
		main_nist_clock_nist_clock_uart_phy_tx_reg <= main_nist_clock_nist_clock_uart_phy_sink_payload_data;
		main_nist_clock_nist_clock_uart_phy_tx_bitcount <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((main_nist_clock_nist_clock_uart_phy_uart_clk_txen & main_nist_clock_nist_clock_uart_phy_tx_busy)) begin
			main_nist_clock_nist_clock_uart_phy_tx_bitcount <= (main_nist_clock_nist_clock_uart_phy_tx_bitcount + 1'd1);
			if ((main_nist_clock_nist_clock_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((main_nist_clock_nist_clock_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					main_nist_clock_nist_clock_uart_phy_tx_busy <= 1'd0;
					main_nist_clock_nist_clock_uart_phy_sink_ack <= 1'd1;
				end else begin
					serial_tx <= main_nist_clock_nist_clock_uart_phy_tx_reg[0];
					main_nist_clock_nist_clock_uart_phy_tx_reg <= {1'd0, main_nist_clock_nist_clock_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (main_nist_clock_nist_clock_uart_phy_tx_busy) begin
		{main_nist_clock_nist_clock_uart_phy_uart_clk_txen, main_nist_clock_nist_clock_uart_phy_phase_accumulator_tx} <= (main_nist_clock_nist_clock_uart_phy_phase_accumulator_tx + main_nist_clock_nist_clock_uart_phy_storage);
	end else begin
		{main_nist_clock_nist_clock_uart_phy_uart_clk_txen, main_nist_clock_nist_clock_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	main_nist_clock_nist_clock_uart_phy_source_stb <= 1'd0;
	main_nist_clock_nist_clock_uart_phy_rx_r <= main_nist_clock_nist_clock_uart_phy_rx;
	if ((~main_nist_clock_nist_clock_uart_phy_rx_busy)) begin
		if (((~main_nist_clock_nist_clock_uart_phy_rx) & main_nist_clock_nist_clock_uart_phy_rx_r)) begin
			main_nist_clock_nist_clock_uart_phy_rx_busy <= 1'd1;
			main_nist_clock_nist_clock_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (main_nist_clock_nist_clock_uart_phy_uart_clk_rxen) begin
			main_nist_clock_nist_clock_uart_phy_rx_bitcount <= (main_nist_clock_nist_clock_uart_phy_rx_bitcount + 1'd1);
			if ((main_nist_clock_nist_clock_uart_phy_rx_bitcount == 1'd0)) begin
				if (main_nist_clock_nist_clock_uart_phy_rx) begin
					main_nist_clock_nist_clock_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((main_nist_clock_nist_clock_uart_phy_rx_bitcount == 4'd9)) begin
					main_nist_clock_nist_clock_uart_phy_rx_busy <= 1'd0;
					if (main_nist_clock_nist_clock_uart_phy_rx) begin
						main_nist_clock_nist_clock_uart_phy_source_payload_data <= main_nist_clock_nist_clock_uart_phy_rx_reg;
						main_nist_clock_nist_clock_uart_phy_source_stb <= 1'd1;
					end
				end else begin
					main_nist_clock_nist_clock_uart_phy_rx_reg <= {main_nist_clock_nist_clock_uart_phy_rx, main_nist_clock_nist_clock_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (main_nist_clock_nist_clock_uart_phy_rx_busy) begin
		{main_nist_clock_nist_clock_uart_phy_uart_clk_rxen, main_nist_clock_nist_clock_uart_phy_phase_accumulator_rx} <= (main_nist_clock_nist_clock_uart_phy_phase_accumulator_rx + main_nist_clock_nist_clock_uart_phy_storage);
	end else begin
		{main_nist_clock_nist_clock_uart_phy_uart_clk_rxen, main_nist_clock_nist_clock_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if (main_nist_clock_nist_clock_uart_tx_clear) begin
		main_nist_clock_nist_clock_uart_tx_pending <= 1'd0;
	end
	main_nist_clock_nist_clock_uart_tx_old_trigger <= main_nist_clock_nist_clock_uart_tx_trigger;
	if (((~main_nist_clock_nist_clock_uart_tx_trigger) & main_nist_clock_nist_clock_uart_tx_old_trigger)) begin
		main_nist_clock_nist_clock_uart_tx_pending <= 1'd1;
	end
	if (main_nist_clock_nist_clock_uart_rx_clear) begin
		main_nist_clock_nist_clock_uart_rx_pending <= 1'd0;
	end
	main_nist_clock_nist_clock_uart_rx_old_trigger <= main_nist_clock_nist_clock_uart_rx_trigger;
	if (((~main_nist_clock_nist_clock_uart_rx_trigger) & main_nist_clock_nist_clock_uart_rx_old_trigger)) begin
		main_nist_clock_nist_clock_uart_rx_pending <= 1'd1;
	end
	if (((main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_we & main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable) & (~main_nist_clock_nist_clock_uart_tx_fifo_replace))) begin
		main_nist_clock_nist_clock_uart_tx_fifo_produce <= (main_nist_clock_nist_clock_uart_tx_fifo_produce + 1'd1);
	end
	if (main_nist_clock_nist_clock_uart_tx_fifo_do_read) begin
		main_nist_clock_nist_clock_uart_tx_fifo_consume <= (main_nist_clock_nist_clock_uart_tx_fifo_consume + 1'd1);
	end
	if (((main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_we & main_nist_clock_nist_clock_uart_tx_fifo_syncfifo_writable) & (~main_nist_clock_nist_clock_uart_tx_fifo_replace))) begin
		if ((~main_nist_clock_nist_clock_uart_tx_fifo_do_read)) begin
			main_nist_clock_nist_clock_uart_tx_fifo_level <= (main_nist_clock_nist_clock_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (main_nist_clock_nist_clock_uart_tx_fifo_do_read) begin
			main_nist_clock_nist_clock_uart_tx_fifo_level <= (main_nist_clock_nist_clock_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_we & main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable) & (~main_nist_clock_nist_clock_uart_rx_fifo_replace))) begin
		main_nist_clock_nist_clock_uart_rx_fifo_produce <= (main_nist_clock_nist_clock_uart_rx_fifo_produce + 1'd1);
	end
	if (main_nist_clock_nist_clock_uart_rx_fifo_do_read) begin
		main_nist_clock_nist_clock_uart_rx_fifo_consume <= (main_nist_clock_nist_clock_uart_rx_fifo_consume + 1'd1);
	end
	if (((main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_we & main_nist_clock_nist_clock_uart_rx_fifo_syncfifo_writable) & (~main_nist_clock_nist_clock_uart_rx_fifo_replace))) begin
		if ((~main_nist_clock_nist_clock_uart_rx_fifo_do_read)) begin
			main_nist_clock_nist_clock_uart_rx_fifo_level <= (main_nist_clock_nist_clock_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (main_nist_clock_nist_clock_uart_rx_fifo_do_read) begin
			main_nist_clock_nist_clock_uart_rx_fifo_level <= (main_nist_clock_nist_clock_uart_rx_fifo_level - 1'd1);
		end
	end
	if (main_nist_clock_nist_clock_timer0_en_storage) begin
		if ((main_nist_clock_nist_clock_timer0_value == 1'd0)) begin
			main_nist_clock_nist_clock_timer0_value <= main_nist_clock_nist_clock_timer0_reload_storage;
		end else begin
			main_nist_clock_nist_clock_timer0_value <= (main_nist_clock_nist_clock_timer0_value - 1'd1);
		end
	end else begin
		main_nist_clock_nist_clock_timer0_value <= main_nist_clock_nist_clock_timer0_load_storage;
	end
	if (main_nist_clock_nist_clock_timer0_update_value_re) begin
		main_nist_clock_nist_clock_timer0_value_status <= main_nist_clock_nist_clock_timer0_value;
	end
	if (main_nist_clock_nist_clock_timer0_zero_clear) begin
		main_nist_clock_nist_clock_timer0_zero_pending <= 1'd0;
	end
	main_nist_clock_nist_clock_timer0_zero_old_trigger <= main_nist_clock_nist_clock_timer0_zero_trigger;
	if (((~main_nist_clock_nist_clock_timer0_zero_trigger) & main_nist_clock_nist_clock_timer0_zero_old_trigger)) begin
		main_nist_clock_nist_clock_timer0_zero_pending <= 1'd1;
	end
	main_nist_clock_ddrphy_n_rddata_en0 <= main_nist_clock_ddrphy_dfi_p0_rddata_en;
	main_nist_clock_ddrphy_n_rddata_en1 <= main_nist_clock_ddrphy_n_rddata_en0;
	main_nist_clock_ddrphy_n_rddata_en2 <= main_nist_clock_ddrphy_n_rddata_en1;
	main_nist_clock_ddrphy_n_rddata_en3 <= main_nist_clock_ddrphy_n_rddata_en2;
	main_nist_clock_ddrphy_n_rddata_en4 <= main_nist_clock_ddrphy_n_rddata_en3;
	main_nist_clock_ddrphy_dfi_p0_rddata_valid <= (main_nist_clock_ddrphy_n_rddata_en4 | main_nist_clock_ddrphy_wlevel_en_storage);
	main_nist_clock_ddrphy_dfi_p1_rddata_valid <= (main_nist_clock_ddrphy_n_rddata_en4 | main_nist_clock_ddrphy_wlevel_en_storage);
	main_nist_clock_ddrphy_dfi_p2_rddata_valid <= (main_nist_clock_ddrphy_n_rddata_en4 | main_nist_clock_ddrphy_wlevel_en_storage);
	main_nist_clock_ddrphy_dfi_p3_rddata_valid <= (main_nist_clock_ddrphy_n_rddata_en4 | main_nist_clock_ddrphy_wlevel_en_storage);
	main_nist_clock_ddrphy_last_wrdata_en <= {main_nist_clock_ddrphy_last_wrdata_en[2:0], main_nist_clock_ddrphy_dfi_p2_wrdata_en};
	if (main_nist_clock_ddrphy_wlevel_en_storage) begin
		main_nist_clock_ddrphy_oe_dqs <= 1'd1;
		main_nist_clock_ddrphy_oe_dq <= 1'd0;
	end else begin
		main_nist_clock_ddrphy_oe_dqs <= main_nist_clock_ddrphy_oe;
		main_nist_clock_ddrphy_oe_dq <= main_nist_clock_ddrphy_oe;
	end
	if (main_nist_clock_nist_clock_inti_p0_rddata_valid) begin
		main_nist_clock_nist_clock_phaseinjector0_status <= main_nist_clock_nist_clock_inti_p0_rddata;
	end
	if (main_nist_clock_nist_clock_inti_p1_rddata_valid) begin
		main_nist_clock_nist_clock_phaseinjector1_status <= main_nist_clock_nist_clock_inti_p1_rddata;
	end
	if (main_nist_clock_nist_clock_inti_p2_rddata_valid) begin
		main_nist_clock_nist_clock_phaseinjector2_status <= main_nist_clock_nist_clock_inti_p2_rddata;
	end
	if (main_nist_clock_nist_clock_inti_p3_rddata_valid) begin
		main_nist_clock_nist_clock_phaseinjector3_status <= main_nist_clock_nist_clock_inti_p3_rddata;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce0) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank0_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank0_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank0_row1 <= main_nist_clock_nist_clock_sdram_controller_bank0_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset0) begin
		main_nist_clock_nist_clock_sdram_controller_bank0_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank0_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce1) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank1_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank1_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank1_row1 <= main_nist_clock_nist_clock_sdram_controller_bank1_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset1) begin
		main_nist_clock_nist_clock_sdram_controller_bank1_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank1_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce2) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank2_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank2_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank2_row1 <= main_nist_clock_nist_clock_sdram_controller_bank2_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset2) begin
		main_nist_clock_nist_clock_sdram_controller_bank2_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank2_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce3) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank3_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank3_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank3_row1 <= main_nist_clock_nist_clock_sdram_controller_bank3_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset3) begin
		main_nist_clock_nist_clock_sdram_controller_bank3_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank3_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce4) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank4_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank4_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank4_row1 <= main_nist_clock_nist_clock_sdram_controller_bank4_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset4) begin
		main_nist_clock_nist_clock_sdram_controller_bank4_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank4_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce5) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank5_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank5_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank5_row1 <= main_nist_clock_nist_clock_sdram_controller_bank5_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset5) begin
		main_nist_clock_nist_clock_sdram_controller_bank5_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank5_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce6) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank6_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank6_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank6_row1 <= main_nist_clock_nist_clock_sdram_controller_bank6_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset6) begin
		main_nist_clock_nist_clock_sdram_controller_bank6_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank6_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_ce7) begin
		if (main_nist_clock_nist_clock_sdram_controller_bank7_open) begin
			main_nist_clock_nist_clock_sdram_controller_bank7_idle <= 1'd0;
			main_nist_clock_nist_clock_sdram_controller_bank7_row1 <= main_nist_clock_nist_clock_sdram_controller_bank7_row0;
		end
	end
	if (main_nist_clock_nist_clock_sdram_controller_reset7) begin
		main_nist_clock_nist_clock_sdram_controller_bank7_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank7_row1 <= 14'd0;
	end
	if (main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_wait) begin
		if ((~main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_done)) begin
			main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count <= (main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count - 1'd1);
		end
	end else begin
		main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count <= 3'd4;
	end
	if (main_nist_clock_nist_clock_sdram_controller_refresh_timer_wait) begin
		if ((~main_nist_clock_nist_clock_sdram_controller_refresh_timer_done)) begin
			main_nist_clock_nist_clock_sdram_controller_refresh_timer_count <= (main_nist_clock_nist_clock_sdram_controller_refresh_timer_count - 1'd1);
		end
	end else begin
		main_nist_clock_nist_clock_sdram_controller_refresh_timer_count <= 10'd975;
	end
	builder_minicon_state <= builder_minicon_next_state;
	main_nist_clock_nist_clock_adr_offset_r <= main_nist_clock_nist_clock_cpulevel_sdram_if_arbitrated_adr[3:0];
	builder_fullmemorywe_state <= builder_fullmemorywe_next_state;
	if ((main_nist_clock_spiflash_i1 == 1'd0)) begin
		main_nist_clock_spiflash_clk <= 1'd1;
		main_nist_clock_spiflash_dqi <= main_nist_clock_spiflash_i0;
	end
	if ((main_nist_clock_spiflash_i1 == 1'd1)) begin
		main_nist_clock_spiflash_i1 <= 1'd0;
		main_nist_clock_spiflash_clk <= 1'd0;
		main_nist_clock_spiflash_sr <= {main_nist_clock_spiflash_sr[27:0], main_nist_clock_spiflash_dqi};
	end else begin
		main_nist_clock_spiflash_i1 <= (main_nist_clock_spiflash_i1 + 1'd1);
	end
	if ((((main_nist_clock_spiflash_bus_cyc & main_nist_clock_spiflash_bus_stb) & (main_nist_clock_spiflash_i1 == 1'd1)) & (main_nist_clock_spiflash_counter == 1'd0))) begin
		main_nist_clock_spiflash_dq_oe <= 1'd1;
		main_nist_clock_spiflash_cs_n1 <= 1'd0;
		main_nist_clock_spiflash_sr[31:0] <= 32'd4294901503;
	end
	if ((main_nist_clock_spiflash_counter == 5'd16)) begin
		main_nist_clock_spiflash_sr[31:8] <= {main_nist_clock_spiflash_bus_adr, {2{1'd0}}};
	end
	if ((main_nist_clock_spiflash_counter == 5'd28)) begin
		main_nist_clock_spiflash_dq_oe <= 1'd0;
	end
	if ((main_nist_clock_spiflash_counter == 7'd66)) begin
		main_nist_clock_spiflash_bus_ack <= 1'd1;
		main_nist_clock_spiflash_cs_n1 <= 1'd1;
	end
	if ((main_nist_clock_spiflash_counter == 7'd67)) begin
		main_nist_clock_spiflash_bus_ack <= 1'd0;
	end
	if ((main_nist_clock_spiflash_counter == 7'd69)) begin
	end
	if ((main_nist_clock_spiflash_counter == 7'd69)) begin
		main_nist_clock_spiflash_counter <= 1'd0;
	end else begin
		if ((main_nist_clock_spiflash_counter != 1'd0)) begin
			main_nist_clock_spiflash_counter <= (main_nist_clock_spiflash_counter + 1'd1);
		end else begin
			if (((main_nist_clock_spiflash_bus_cyc & main_nist_clock_spiflash_bus_stb) & (main_nist_clock_spiflash_i1 == 1'd1))) begin
				main_nist_clock_spiflash_counter <= 1'd1;
			end
		end
	end
	if (main_ethphy_update_mode) begin
		main_ethphy_mode0 <= main_ethphy_mode1;
	end
	if (main_ethphy_sys_counter_reset) begin
		main_ethphy_sys_counter <= 1'd0;
	end else begin
		if (main_ethphy_sys_counter_ce) begin
			main_ethphy_sys_counter <= (main_ethphy_sys_counter + 1'd1);
		end
	end
	main_ethphy_toggle_o_r <= main_ethphy_toggle_o;
	builder_liteethphygmiimii_state <= builder_liteethphygmiimii_next_state;
	if (main_ps_preamble_error_o) begin
		main_preamble_errors_status <= (main_preamble_errors_status + 1'd1);
	end
	if (main_ps_crc_error_o) begin
		main_crc_errors_status <= (main_crc_errors_status + 1'd1);
	end
	main_ps_preamble_error_toggle_o_r <= main_ps_preamble_error_toggle_o;
	main_ps_crc_error_toggle_o_r <= main_ps_crc_error_toggle_o;
	main_tx_cdc_graycounter0_q_binary <= main_tx_cdc_graycounter0_q_next_binary;
	main_tx_cdc_graycounter0_q <= main_tx_cdc_graycounter0_q_next;
	main_rx_cdc_graycounter1_q_binary <= main_rx_cdc_graycounter1_q_next_binary;
	main_rx_cdc_graycounter1_q <= main_rx_cdc_graycounter1_q_next;
	if (main_writer_counter_reset) begin
		main_writer_counter <= 1'd0;
	end else begin
		if (main_writer_counter_ce) begin
			main_writer_counter <= (main_writer_counter + main_writer_increment);
		end
	end
	if (main_writer_slot_ce) begin
		main_writer_slot <= (main_writer_slot + 1'd1);
	end
	if (((main_writer_fifo_syncfifo_we & main_writer_fifo_syncfifo_writable) & (~main_writer_fifo_replace))) begin
		main_writer_fifo_produce <= (main_writer_fifo_produce + 1'd1);
	end
	if (main_writer_fifo_do_read) begin
		main_writer_fifo_consume <= (main_writer_fifo_consume + 1'd1);
	end
	if (((main_writer_fifo_syncfifo_we & main_writer_fifo_syncfifo_writable) & (~main_writer_fifo_replace))) begin
		if ((~main_writer_fifo_do_read)) begin
			main_writer_fifo_level <= (main_writer_fifo_level + 1'd1);
		end
	end else begin
		if (main_writer_fifo_do_read) begin
			main_writer_fifo_level <= (main_writer_fifo_level - 1'd1);
		end
	end
	builder_liteethmacsramwriter_state <= builder_liteethmacsramwriter_next_state;
	if (main_writer_errors_status_next_value_ce) begin
		main_writer_errors_status <= main_writer_errors_status_next_value;
	end
	if (main_reader_counter_reset) begin
		main_reader_counter <= 1'd0;
	end else begin
		if (main_reader_counter_ce) begin
			main_reader_counter <= (main_reader_counter + 3'd4);
		end
	end
	main_reader_last_d <= main_reader_last;
	if (main_reader_done_clear) begin
		main_reader_done_pending <= 1'd0;
	end
	if (main_reader_done_trigger) begin
		main_reader_done_pending <= 1'd1;
	end
	if (((main_reader_fifo_syncfifo_we & main_reader_fifo_syncfifo_writable) & (~main_reader_fifo_replace))) begin
		main_reader_fifo_produce <= (main_reader_fifo_produce + 1'd1);
	end
	if (main_reader_fifo_do_read) begin
		main_reader_fifo_consume <= (main_reader_fifo_consume + 1'd1);
	end
	if (((main_reader_fifo_syncfifo_we & main_reader_fifo_syncfifo_writable) & (~main_reader_fifo_replace))) begin
		if ((~main_reader_fifo_do_read)) begin
			main_reader_fifo_level <= (main_reader_fifo_level + 1'd1);
		end
	end else begin
		if (main_reader_fifo_do_read) begin
			main_reader_fifo_level <= (main_reader_fifo_level - 1'd1);
		end
	end
	builder_liteethmacsramreader_state <= builder_liteethmacsramreader_next_state;
	main_sram0_bus_ack0 <= 1'd0;
	if (((main_sram0_bus_cyc0 & main_sram0_bus_stb0) & (~main_sram0_bus_ack0))) begin
		main_sram0_bus_ack0 <= 1'd1;
	end
	main_sram1_bus_ack0 <= 1'd0;
	if (((main_sram1_bus_cyc0 & main_sram1_bus_stb0) & (~main_sram1_bus_ack0))) begin
		main_sram1_bus_ack0 <= 1'd1;
	end
	main_sram2_bus_ack0 <= 1'd0;
	if (((main_sram2_bus_cyc0 & main_sram2_bus_stb0) & (~main_sram2_bus_ack0))) begin
		main_sram2_bus_ack0 <= 1'd1;
	end
	main_sram3_bus_ack0 <= 1'd0;
	if (((main_sram3_bus_cyc0 & main_sram3_bus_stb0) & (~main_sram3_bus_ack0))) begin
		main_sram3_bus_ack0 <= 1'd1;
	end
	main_sram0_bus_ack1 <= 1'd0;
	if (((main_sram0_bus_cyc1 & main_sram0_bus_stb1) & (~main_sram0_bus_ack1))) begin
		main_sram0_bus_ack1 <= 1'd1;
	end
	main_sram1_bus_ack1 <= 1'd0;
	if (((main_sram1_bus_cyc1 & main_sram1_bus_stb1) & (~main_sram1_bus_ack1))) begin
		main_sram1_bus_ack1 <= 1'd1;
	end
	main_sram2_bus_ack1 <= 1'd0;
	if (((main_sram2_bus_cyc1 & main_sram2_bus_stb1) & (~main_sram2_bus_ack1))) begin
		main_sram2_bus_ack1 <= 1'd1;
	end
	main_sram3_bus_ack1 <= 1'd0;
	if (((main_sram3_bus_cyc1 & main_sram3_bus_stb1) & (~main_sram3_bus_ack1))) begin
		main_sram3_bus_ack1 <= 1'd1;
	end
	main_slave_sel_r <= main_slave_sel;
	case (builder_grant)
		1'd0: begin
			if ((~builder_request[0])) begin
				if (builder_request[1]) begin
					builder_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_request[1])) begin
				if (builder_request[0]) begin
					builder_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_slave_sel_r <= builder_slave_sel;
	main_mailbox_i1_dat_r <= builder_sync_rhs_array_muxed2;
	main_mailbox_i1_ack <= 1'd0;
	if (((main_mailbox_i1_cyc & main_mailbox_i1_stb) & (~main_mailbox_i1_ack))) begin
		main_mailbox_i1_ack <= 1'd1;
		if (main_mailbox_i1_we) begin
			builder_sync_t_t_array_muxed0 = main_mailbox_i1_dat_w;
			case (main_mailbox_i1_adr[1:0])
				1'd0: begin
					main_mailbox0 <= builder_sync_t_t_array_muxed0;
				end
				1'd1: begin
					main_mailbox1 <= builder_sync_t_t_array_muxed0;
				end
				default: begin
					main_mailbox2 <= builder_sync_t_t_array_muxed0;
				end
			endcase
		end
	end
	main_mailbox_i2_dat_r <= builder_sync_rhs_array_muxed3;
	main_mailbox_i2_ack <= 1'd0;
	if (((main_mailbox_i2_cyc & main_mailbox_i2_stb) & (~main_mailbox_i2_ack))) begin
		main_mailbox_i2_ack <= 1'd1;
		if (main_mailbox_i2_we) begin
			builder_sync_t_t_array_muxed1 = main_mailbox_i2_dat_w;
			case (main_mailbox_i2_adr[1:0])
				1'd0: begin
					main_mailbox0 <= builder_sync_t_t_array_muxed1;
				end
				1'd1: begin
					main_mailbox1 <= builder_sync_t_t_array_muxed1;
				end
				default: begin
					main_mailbox2 <= builder_sync_t_t_array_muxed1;
				end
			endcase
		end
	end
	if (main_en_storage) begin
		if ((main_value == 1'd0)) begin
			main_value <= main_reload_storage;
		end else begin
			main_value <= (main_value - 1'd1);
		end
	end else begin
		main_value <= main_load_storage;
	end
	if (main_update_value_re) begin
		main_value_status <= main_value;
	end
	if (main_zero_clear) begin
		main_zero_pending <= 1'd0;
	end
	main_zero_old_trigger <= main_zero_trigger;
	if (((~main_zero_trigger) & main_zero_old_trigger)) begin
		main_zero_pending <= 1'd1;
	end
	main_o <= main_value_sys;
	main_rtio_core_cmd_reset <= main_rtio_core_reset_re;
	main_rtio_core_cmd_reset_phy <= main_rtio_core_reset_phy_re;
	main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= (main_coarse_ts_sys + 5'd16);
	if (main_rtio_core_async_error_re) begin
		if (main_rtio_core_async_error_r[0]) begin
			main_rtio_core_o_collision <= 1'd0;
		end
		if (main_rtio_core_async_error_r[1]) begin
			main_rtio_core_o_busy <= 1'd0;
		end
		if (main_rtio_core_async_error_r[2]) begin
			main_rtio_core_o_sequence_error <= 1'd0;
		end
	end
	if (main_rtio_core_o_collision_sync_o) begin
		main_rtio_core_o_collision <= 1'd1;
		if ((~main_rtio_core_o_collision)) begin
			main_rtio_core_collision_channel_status <= main_rtio_core_o_collision_sync_data_o;
		end
	end
	if (main_rtio_core_o_busy_sync_o) begin
		main_rtio_core_o_busy <= 1'd1;
		if ((~main_rtio_core_o_busy)) begin
			main_rtio_core_busy_channel_status <= main_rtio_core_o_busy_sync_data_o;
		end
	end
	if (main_rtio_core_outputs_lanedistributor_sequence_error) begin
		main_rtio_core_o_sequence_error <= 1'd1;
		if ((~main_rtio_core_o_sequence_error)) begin
			main_rtio_core_sequence_error_channel_status <= main_rtio_core_outputs_lanedistributor_sequence_error_channel;
		end
	end
	if (main_rtio_now_hi_re) begin
		main_rtio_now_hi_backing <= main_rtio_now_hi_r;
	end
	if (main_rtio_now_lo_re) begin
		main_rtio_now <= {main_rtio_now_hi_backing, main_rtio_now_lo_r};
	end
	if (main_rtio_counter_update_re) begin
		main_rtio_counter_status <= main_full_ts_sys;
	end
	case (main_csrbank0_bus_adr[4:0])
		1'd0: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_target0_w;
		end
		1'd1: begin
			main_csrbank0_bus_dat_r <= main_rtio_now_hi_w;
		end
		2'd2: begin
			main_csrbank0_bus_dat_r <= main_rtio_now_lo_w;
		end
		2'd3: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data15_w;
		end
		3'd4: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data14_w;
		end
		3'd5: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data13_w;
		end
		3'd6: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data12_w;
		end
		3'd7: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data11_w;
		end
		4'd8: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data10_w;
		end
		4'd9: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data9_w;
		end
		4'd10: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data8_w;
		end
		4'd11: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data7_w;
		end
		4'd12: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data6_w;
		end
		4'd13: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data5_w;
		end
		4'd14: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data4_w;
		end
		4'd15: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data3_w;
		end
		5'd16: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data2_w;
		end
		5'd17: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data1_w;
		end
		5'd18: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_data0_w;
		end
		5'd19: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_o_status_w;
		end
		5'd20: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_timeout1_w;
		end
		5'd21: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_timeout0_w;
		end
		5'd22: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_data_w;
		end
		5'd23: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_timestamp1_w;
		end
		5'd24: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_timestamp0_w;
		end
		5'd25: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_i_status_w;
		end
		5'd26: begin
			main_csrbank0_bus_dat_r <= main_rtio_i_overflow_reset_w;
		end
		5'd27: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_counter1_w;
		end
		5'd28: begin
			main_csrbank0_bus_dat_r <= main_csrbank0_counter0_w;
		end
		5'd29: begin
			main_csrbank0_bus_dat_r <= main_rtio_counter_update_w;
		end
	endcase
	if (main_csrbank0_bus_ack) begin
		main_csrbank0_bus_ack <= 1'd0;
	end else begin
		if ((main_csrbank0_bus_cyc & main_csrbank0_bus_stb)) begin
			main_csrbank0_bus_ack <= 1'd1;
		end
	end
	if (main_csrbank0_target0_re) begin
		main_rtio_target_storage_full[31:0] <= main_csrbank0_target0_r;
	end
	main_rtio_target_re <= main_csrbank0_target0_re;
	if (main_rtio_o_data_we) begin
		main_rtio_o_data_storage_full <= (main_rtio_o_data_dat_w <<< 1'd0);
	end
	if (main_csrbank0_o_data15_re) begin
		main_rtio_o_data_storage_full[511:480] <= main_csrbank0_o_data15_r;
	end
	if (main_csrbank0_o_data14_re) begin
		main_rtio_o_data_storage_full[479:448] <= main_csrbank0_o_data14_r;
	end
	if (main_csrbank0_o_data13_re) begin
		main_rtio_o_data_storage_full[447:416] <= main_csrbank0_o_data13_r;
	end
	if (main_csrbank0_o_data12_re) begin
		main_rtio_o_data_storage_full[415:384] <= main_csrbank0_o_data12_r;
	end
	if (main_csrbank0_o_data11_re) begin
		main_rtio_o_data_storage_full[383:352] <= main_csrbank0_o_data11_r;
	end
	if (main_csrbank0_o_data10_re) begin
		main_rtio_o_data_storage_full[351:320] <= main_csrbank0_o_data10_r;
	end
	if (main_csrbank0_o_data9_re) begin
		main_rtio_o_data_storage_full[319:288] <= main_csrbank0_o_data9_r;
	end
	if (main_csrbank0_o_data8_re) begin
		main_rtio_o_data_storage_full[287:256] <= main_csrbank0_o_data8_r;
	end
	if (main_csrbank0_o_data7_re) begin
		main_rtio_o_data_storage_full[255:224] <= main_csrbank0_o_data7_r;
	end
	if (main_csrbank0_o_data6_re) begin
		main_rtio_o_data_storage_full[223:192] <= main_csrbank0_o_data6_r;
	end
	if (main_csrbank0_o_data5_re) begin
		main_rtio_o_data_storage_full[191:160] <= main_csrbank0_o_data5_r;
	end
	if (main_csrbank0_o_data4_re) begin
		main_rtio_o_data_storage_full[159:128] <= main_csrbank0_o_data4_r;
	end
	if (main_csrbank0_o_data3_re) begin
		main_rtio_o_data_storage_full[127:96] <= main_csrbank0_o_data3_r;
	end
	if (main_csrbank0_o_data2_re) begin
		main_rtio_o_data_storage_full[95:64] <= main_csrbank0_o_data2_r;
	end
	if (main_csrbank0_o_data1_re) begin
		main_rtio_o_data_storage_full[63:32] <= main_csrbank0_o_data1_r;
	end
	if (main_csrbank0_o_data0_re) begin
		main_rtio_o_data_storage_full[31:0] <= main_csrbank0_o_data0_r;
	end
	main_rtio_o_data_re <= main_csrbank0_o_data0_re;
	if (main_csrbank0_i_timeout1_re) begin
		main_rtio_i_timeout_storage_full[63:32] <= main_csrbank0_i_timeout1_r;
	end
	if (main_csrbank0_i_timeout0_re) begin
		main_rtio_i_timeout_storage_full[31:0] <= main_csrbank0_i_timeout0_r;
	end
	main_rtio_i_timeout_re <= main_csrbank0_i_timeout0_re;
	case (main_csrbank1_bus_adr[3:0])
		1'd0: begin
			main_csrbank1_bus_dat_r <= main_dma_enable_enable_w;
		end
		1'd1: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_base_address1_w;
		end
		2'd2: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_base_address0_w;
		end
		2'd3: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_time_offset1_w;
		end
		3'd4: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_time_offset0_w;
		end
		3'd5: begin
			main_csrbank1_bus_dat_r <= main_dma_cri_master_error_w;
		end
		3'd6: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_error_channel_w;
		end
		3'd7: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_error_timestamp1_w;
		end
		4'd8: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_error_timestamp0_w;
		end
		4'd9: begin
			main_csrbank1_bus_dat_r <= main_csrbank1_error_address_w;
		end
	endcase
	if (main_csrbank1_bus_ack) begin
		main_csrbank1_bus_ack <= 1'd0;
	end else begin
		if ((main_csrbank1_bus_cyc & main_csrbank1_bus_stb)) begin
			main_csrbank1_bus_ack <= 1'd1;
		end
	end
	if (main_csrbank1_base_address1_re) begin
		main_dma_dma_storage_full[35:32] <= main_csrbank1_base_address1_r;
	end
	if (main_csrbank1_base_address0_re) begin
		main_dma_dma_storage_full[31:0] <= main_csrbank1_base_address0_r;
	end
	main_dma_dma_re <= main_csrbank1_base_address0_re;
	if (main_csrbank1_time_offset1_re) begin
		main_dma_time_offset_storage_full[63:32] <= main_csrbank1_time_offset1_r;
	end
	if (main_csrbank1_time_offset0_re) begin
		main_dma_time_offset_storage_full[31:0] <= main_csrbank1_time_offset0_r;
	end
	main_dma_time_offset_re <= main_csrbank1_time_offset0_re;
	main_cri_con_selected <= main_cri_con_shared_chan_sel[23:16];
	case (main_csrbank2_bus_adr[0])
		1'd0: begin
			main_csrbank2_bus_dat_r <= main_csrbank2_selected0_w;
		end
	endcase
	if (main_csrbank2_bus_ack) begin
		main_csrbank2_bus_ack <= 1'd0;
	end else begin
		if ((main_csrbank2_bus_cyc & main_csrbank2_bus_stb)) begin
			main_csrbank2_bus_ack <= 1'd1;
		end
	end
	if (main_csrbank2_selected0_re) begin
		main_cri_con_storage_full[1:0] <= main_csrbank2_selected0_r;
	end
	main_cri_con_re <= main_csrbank2_selected0_re;
	if (main_mon_value_update_re) begin
		main_mon_status <= builder_sync_t_rhs_array_muxed2;
	end
	main_mon_bussynchronizer28_ping_o1 <= main_mon_bussynchronizer28_ping_o0;
	if (main_mon_bussynchronizer28_ping_o1) begin
		main_mon_bussynchronizer28_o <= main_mon_bussynchronizer28_obuffer;
	end
	main_mon_bussynchronizer28_ping_toggle_o_r <= main_mon_bussynchronizer28_ping_toggle_o;
	if (main_mon_bussynchronizer28_pong_i) begin
		main_mon_bussynchronizer28_pong_toggle_i <= (~main_mon_bussynchronizer28_pong_toggle_i);
	end
	main_mon_bussynchronizer29_ping_o1 <= main_mon_bussynchronizer29_ping_o0;
	if (main_mon_bussynchronizer29_ping_o1) begin
		main_mon_bussynchronizer29_o <= main_mon_bussynchronizer29_obuffer;
	end
	main_mon_bussynchronizer29_ping_toggle_o_r <= main_mon_bussynchronizer29_ping_toggle_o;
	if (main_mon_bussynchronizer29_pong_i) begin
		main_mon_bussynchronizer29_pong_toggle_i <= (~main_mon_bussynchronizer29_pong_toggle_i);
	end
	main_mon_bussynchronizer30_ping_o1 <= main_mon_bussynchronizer30_ping_o0;
	if (main_mon_bussynchronizer30_ping_o1) begin
		main_mon_bussynchronizer30_o <= main_mon_bussynchronizer30_obuffer;
	end
	main_mon_bussynchronizer30_ping_toggle_o_r <= main_mon_bussynchronizer30_ping_toggle_o;
	if (main_mon_bussynchronizer30_pong_i) begin
		main_mon_bussynchronizer30_pong_toggle_i <= (~main_mon_bussynchronizer30_pong_toggle_i);
	end
	main_mon_bussynchronizer31_ping_o1 <= main_mon_bussynchronizer31_ping_o0;
	if (main_mon_bussynchronizer31_ping_o1) begin
		main_mon_bussynchronizer31_o <= main_mon_bussynchronizer31_obuffer;
	end
	main_mon_bussynchronizer31_ping_toggle_o_r <= main_mon_bussynchronizer31_ping_toggle_o;
	if (main_mon_bussynchronizer31_pong_i) begin
		main_mon_bussynchronizer31_pong_toggle_i <= (~main_mon_bussynchronizer31_pong_toggle_i);
	end
	main_mon_bussynchronizer32_ping_o1 <= main_mon_bussynchronizer32_ping_o0;
	if (main_mon_bussynchronizer32_ping_o1) begin
		main_mon_bussynchronizer32_o <= main_mon_bussynchronizer32_obuffer;
	end
	main_mon_bussynchronizer32_ping_toggle_o_r <= main_mon_bussynchronizer32_ping_toggle_o;
	if (main_mon_bussynchronizer32_pong_i) begin
		main_mon_bussynchronizer32_pong_toggle_i <= (~main_mon_bussynchronizer32_pong_toggle_i);
	end
	main_mon_bussynchronizer33_ping_o1 <= main_mon_bussynchronizer33_ping_o0;
	if (main_mon_bussynchronizer33_ping_o1) begin
		main_mon_bussynchronizer33_o <= main_mon_bussynchronizer33_obuffer;
	end
	main_mon_bussynchronizer33_ping_toggle_o_r <= main_mon_bussynchronizer33_ping_toggle_o;
	if (main_mon_bussynchronizer33_pong_i) begin
		main_mon_bussynchronizer33_pong_toggle_i <= (~main_mon_bussynchronizer33_pong_toggle_i);
	end
	main_mon_bussynchronizer34_ping_o1 <= main_mon_bussynchronizer34_ping_o0;
	if (main_mon_bussynchronizer34_ping_o1) begin
		main_mon_bussynchronizer34_o <= main_mon_bussynchronizer34_obuffer;
	end
	main_mon_bussynchronizer34_ping_toggle_o_r <= main_mon_bussynchronizer34_ping_toggle_o;
	if (main_mon_bussynchronizer34_pong_i) begin
		main_mon_bussynchronizer34_pong_toggle_i <= (~main_mon_bussynchronizer34_pong_toggle_i);
	end
	main_mon_bussynchronizer35_ping_o1 <= main_mon_bussynchronizer35_ping_o0;
	if (main_mon_bussynchronizer35_ping_o1) begin
		main_mon_bussynchronizer35_o <= main_mon_bussynchronizer35_obuffer;
	end
	main_mon_bussynchronizer35_ping_toggle_o_r <= main_mon_bussynchronizer35_ping_toggle_o;
	if (main_mon_bussynchronizer35_pong_i) begin
		main_mon_bussynchronizer35_pong_toggle_i <= (~main_mon_bussynchronizer35_pong_toggle_i);
	end
	main_mon_bussynchronizer36_ping_o1 <= main_mon_bussynchronizer36_ping_o0;
	if (main_mon_bussynchronizer36_ping_o1) begin
		main_mon_bussynchronizer36_o <= main_mon_bussynchronizer36_obuffer;
	end
	main_mon_bussynchronizer36_ping_toggle_o_r <= main_mon_bussynchronizer36_ping_toggle_o;
	if (main_mon_bussynchronizer36_pong_i) begin
		main_mon_bussynchronizer36_pong_toggle_i <= (~main_mon_bussynchronizer36_pong_toggle_i);
	end
	main_mon_bussynchronizer37_ping_o1 <= main_mon_bussynchronizer37_ping_o0;
	if (main_mon_bussynchronizer37_ping_o1) begin
		main_mon_bussynchronizer37_o <= main_mon_bussynchronizer37_obuffer;
	end
	main_mon_bussynchronizer37_ping_toggle_o_r <= main_mon_bussynchronizer37_ping_toggle_o;
	if (main_mon_bussynchronizer37_pong_i) begin
		main_mon_bussynchronizer37_pong_toggle_i <= (~main_mon_bussynchronizer37_pong_toggle_i);
	end
	main_mon_bussynchronizer38_ping_o1 <= main_mon_bussynchronizer38_ping_o0;
	if (main_mon_bussynchronizer38_ping_o1) begin
		main_mon_bussynchronizer38_o <= main_mon_bussynchronizer38_obuffer;
	end
	main_mon_bussynchronizer38_ping_toggle_o_r <= main_mon_bussynchronizer38_ping_toggle_o;
	if (main_mon_bussynchronizer38_pong_i) begin
		main_mon_bussynchronizer38_pong_toggle_i <= (~main_mon_bussynchronizer38_pong_toggle_i);
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd0)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys0 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd0)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys1 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd1)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys2 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 1'd1)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys3 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd2)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys4 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd2)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys5 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys6 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys7 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 2'd3)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys8 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd4)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys9 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd4)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys10 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd5)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys11 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd5)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys12 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd6)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys13 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd6)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys14 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys15 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys16 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 3'd7)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys17 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd8)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys18 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd8)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys19 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd9)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys20 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd9)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys21 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd10)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys22 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd10)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys23 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd11)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys24 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd11)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys25 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd11)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys26 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd12)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys27 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd12)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys28 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd13)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys29 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd13)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys30 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd14)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys31 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd14)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys32 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd15)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys33 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd15)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys34 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 4'd15)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys35 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd16)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys36 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd16)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys37 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd16)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys38 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd17)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys39 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd17)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys40 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd17)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys41 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd18)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys42 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd18)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys43 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd18)) & (main_inj_override_sel_storage == 2'd2))) begin
		main_inj_o_sys44 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd19)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys45 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd19)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys46 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd20)) & (main_inj_override_sel_storage == 1'd0))) begin
		main_inj_o_sys47 <= main_inj_value_r;
	end
	if (((main_inj_value_re & (main_inj_chan_sel_storage == 5'd20)) & (main_inj_override_sel_storage == 1'd1))) begin
		main_inj_o_sys48 <= main_inj_value_r;
	end
	main_rtio_analyzer_enable_r <= main_rtio_analyzer_enable_storage;
	if ((main_rtio_analyzer_enable_storage & (~main_rtio_analyzer_enable_r))) begin
		main_rtio_analyzer_busy_status <= 1'd1;
	end
	if (((main_rtio_analyzer_dma_sink_stb & main_rtio_analyzer_dma_sink_ack) & main_rtio_analyzer_dma_sink_eop)) begin
		main_rtio_analyzer_busy_status <= 1'd0;
	end
	main_rtio_analyzer_message_encoder_read_wait_event_r <= main_rtio_core_cri_i_status[2];
	main_rtio_analyzer_message_encoder_just_written <= (main_rtio_core_cri_cmd == 1'd1);
	main_rtio_analyzer_message_encoder_enable_r <= main_rtio_analyzer_enable_storage;
	if (((~main_rtio_analyzer_enable_storage) & main_rtio_analyzer_message_encoder_enable_r)) begin
		main_rtio_analyzer_message_encoder_stopping <= 1'd1;
	end
	if ((~main_rtio_analyzer_message_encoder_stopping)) begin
		if (main_rtio_analyzer_message_encoder_exception_stb) begin
			main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_exception_padding1, main_rtio_analyzer_message_encoder_exception_exception_type, main_rtio_analyzer_message_encoder_exception_rtio_counter, main_rtio_analyzer_message_encoder_exception_padding0, main_rtio_analyzer_message_encoder_exception_channel, main_rtio_analyzer_message_encoder_exception_message_type};
		end else begin
			main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_input_output_data, main_rtio_analyzer_message_encoder_input_output_address_padding, main_rtio_analyzer_message_encoder_input_output_rtio_counter, main_rtio_analyzer_message_encoder_input_output_timestamp, main_rtio_analyzer_message_encoder_input_output_channel, main_rtio_analyzer_message_encoder_input_output_message_type};
		end
		main_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_rtio_analyzer_message_encoder_source_stb <= (main_rtio_analyzer_enable_storage & (main_rtio_analyzer_message_encoder_input_output_stb | main_rtio_analyzer_message_encoder_exception_stb));
		if (main_rtio_analyzer_message_encoder_overflow_reset_re) begin
			main_rtio_analyzer_message_encoder_status <= 1'd0;
		end
		if ((main_rtio_analyzer_message_encoder_source_stb & (~main_rtio_analyzer_message_encoder_source_ack))) begin
			main_rtio_analyzer_message_encoder_status <= 1'd1;
		end
	end else begin
		main_rtio_analyzer_message_encoder_source_payload_data <= {main_rtio_analyzer_message_encoder_stopped_padding1, main_rtio_analyzer_message_encoder_stopped_rtio_counter, main_rtio_analyzer_message_encoder_stopped_padding0, main_rtio_analyzer_message_encoder_stopped_message_type};
		main_rtio_analyzer_message_encoder_source_eop <= 1'd1;
		main_rtio_analyzer_message_encoder_source_stb <= 1'd1;
		if (main_rtio_analyzer_message_encoder_source_ack) begin
			main_rtio_analyzer_message_encoder_stopping <= 1'd0;
		end
	end
	if (main_rtio_analyzer_fifo_syncfifo_re) begin
		main_rtio_analyzer_fifo_readable <= 1'd1;
	end else begin
		if (main_rtio_analyzer_fifo_re) begin
			main_rtio_analyzer_fifo_readable <= 1'd0;
		end
	end
	if (((main_rtio_analyzer_fifo_syncfifo_we & main_rtio_analyzer_fifo_syncfifo_writable) & (~main_rtio_analyzer_fifo_replace))) begin
		main_rtio_analyzer_fifo_produce <= (main_rtio_analyzer_fifo_produce + 1'd1);
	end
	if (main_rtio_analyzer_fifo_do_read) begin
		main_rtio_analyzer_fifo_consume <= (main_rtio_analyzer_fifo_consume + 1'd1);
	end
	if (((main_rtio_analyzer_fifo_syncfifo_we & main_rtio_analyzer_fifo_syncfifo_writable) & (~main_rtio_analyzer_fifo_replace))) begin
		if ((~main_rtio_analyzer_fifo_do_read)) begin
			main_rtio_analyzer_fifo_level0 <= (main_rtio_analyzer_fifo_level0 + 1'd1);
		end
	end else begin
		if (main_rtio_analyzer_fifo_do_read) begin
			main_rtio_analyzer_fifo_level0 <= (main_rtio_analyzer_fifo_level0 - 1'd1);
		end
	end
	if (main_rtio_analyzer_converter_source_ack) begin
		main_rtio_analyzer_converter_strobe_all <= 1'd0;
	end
	if (main_rtio_analyzer_converter_load_part) begin
		if (((main_rtio_analyzer_converter_demux == 1'd1) | main_rtio_analyzer_converter_sink_eop)) begin
			main_rtio_analyzer_converter_demux <= 1'd0;
			main_rtio_analyzer_converter_strobe_all <= 1'd1;
		end else begin
			main_rtio_analyzer_converter_demux <= (main_rtio_analyzer_converter_demux + 1'd1);
		end
	end
	if ((main_rtio_analyzer_converter_source_stb & main_rtio_analyzer_converter_source_ack)) begin
		main_rtio_analyzer_converter_source_eop <= main_rtio_analyzer_converter_sink_eop;
	end else begin
		if ((main_rtio_analyzer_converter_sink_stb & main_rtio_analyzer_converter_sink_ack)) begin
			main_rtio_analyzer_converter_source_eop <= (main_rtio_analyzer_converter_sink_eop | main_rtio_analyzer_converter_source_eop);
		end
	end
	if (main_rtio_analyzer_converter_load_part) begin
		case (main_rtio_analyzer_converter_demux)
			1'd0: begin
				main_rtio_analyzer_converter_source_payload_data[511:256] <= main_rtio_analyzer_converter_sink_payload_data;
			end
			1'd1: begin
				main_rtio_analyzer_converter_source_payload_data[255:0] <= main_rtio_analyzer_converter_sink_payload_data;
			end
		endcase
	end
	if (main_rtio_analyzer_converter_load_part) begin
		main_rtio_analyzer_converter_source_payload_valid_token_count <= (main_rtio_analyzer_converter_demux + 1'd1);
	end
	if (main_rtio_analyzer_dma_reset_re) begin
		main_interface1_bus_adr <= main_rtio_analyzer_dma_base_address_storage;
	end
	if (main_interface1_bus_ack) begin
		if ((main_interface1_bus_adr == main_rtio_analyzer_dma_last_address_storage)) begin
			main_interface1_bus_adr <= main_rtio_analyzer_dma_base_address_storage;
		end else begin
			main_interface1_bus_adr <= (main_interface1_bus_adr + 1'd1);
		end
	end
	if (main_rtio_analyzer_dma_reset_re) begin
		main_rtio_analyzer_dma_message_count <= 1'd0;
	end
	if (main_interface1_bus_ack) begin
		main_rtio_analyzer_dma_message_count <= (main_rtio_analyzer_dma_message_count + main_rtio_analyzer_dma_sink_payload_valid_token_count);
	end
	case (builder_sdram_cpulevel_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_cpulevel_arbiter_request[0])) begin
				if (builder_sdram_cpulevel_arbiter_request[1]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_cpulevel_arbiter_request[1])) begin
				if (builder_sdram_cpulevel_arbiter_request[0]) begin
					builder_sdram_cpulevel_arbiter_grant <= 1'd0;
				end
			end
		end
	endcase
	case (builder_sdram_native_arbiter_grant)
		1'd0: begin
			if ((~builder_sdram_native_arbiter_request[0])) begin
				if (builder_sdram_native_arbiter_request[1]) begin
					builder_sdram_native_arbiter_grant <= 1'd1;
				end else begin
					if (builder_sdram_native_arbiter_request[2]) begin
						builder_sdram_native_arbiter_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~builder_sdram_native_arbiter_request[1])) begin
				if (builder_sdram_native_arbiter_request[2]) begin
					builder_sdram_native_arbiter_grant <= 2'd2;
				end else begin
					if (builder_sdram_native_arbiter_request[0]) begin
						builder_sdram_native_arbiter_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~builder_sdram_native_arbiter_request[2])) begin
				if (builder_sdram_native_arbiter_request[0]) begin
					builder_sdram_native_arbiter_grant <= 1'd0;
				end else begin
					if (builder_sdram_native_arbiter_request[1]) begin
						builder_sdram_native_arbiter_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	case (builder_nist_clock_grant)
		1'd0: begin
			if ((~builder_nist_clock_request[0])) begin
				if (builder_nist_clock_request[1]) begin
					builder_nist_clock_grant <= 1'd1;
				end
			end
		end
		1'd1: begin
			if ((~builder_nist_clock_request[1])) begin
				if (builder_nist_clock_request[0]) begin
					builder_nist_clock_grant <= 1'd0;
				end
			end
		end
	endcase
	builder_nist_clock_slave_sel_r <= builder_nist_clock_slave_sel;
	builder_nist_clock_interface0_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank0_sel) begin
		case (builder_nist_clock_interface0_bank_bus_adr[3:0])
			1'd0: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= builder_nist_clock_csrbank0_wlevel_en0_w;
			end
			1'd1: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_wlevel_strobe_w;
			end
			2'd2: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= builder_nist_clock_csrbank0_dly_sel0_w;
			end
			2'd3: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_rdly_dq_rst_w;
			end
			3'd4: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_rdly_dq_inc_w;
			end
			3'd5: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_rdly_dq_bitslip_w;
			end
			3'd6: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_wdly_dq_rst_w;
			end
			3'd7: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_wdly_dq_inc_w;
			end
			4'd8: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_wdly_dqs_rst_w;
			end
			4'd9: begin
				builder_nist_clock_interface0_bank_bus_dat_r <= main_nist_clock_ddrphy_wdly_dqs_inc_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank0_wlevel_en0_re) begin
		main_nist_clock_ddrphy_wlevel_en_storage_full <= builder_nist_clock_csrbank0_wlevel_en0_r;
	end
	main_nist_clock_ddrphy_wlevel_en_re <= builder_nist_clock_csrbank0_wlevel_en0_re;
	if (builder_nist_clock_csrbank0_dly_sel0_re) begin
		main_nist_clock_ddrphy_dly_sel_storage_full[7:0] <= builder_nist_clock_csrbank0_dly_sel0_r;
	end
	main_nist_clock_ddrphy_dly_sel_re <= builder_nist_clock_csrbank0_dly_sel0_re;
	builder_nist_clock_interface1_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank1_sel) begin
		case (builder_nist_clock_interface1_bank_bus_adr[7:0])
			1'd0: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_control0_w;
			end
			1'd1: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_command0_w;
			end
			2'd2: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= main_nist_clock_nist_clock_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_address1_w;
			end
			3'd4: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_address0_w;
			end
			3'd5: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_baddress0_w;
			end
			3'd6: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata15_w;
			end
			3'd7: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata14_w;
			end
			4'd8: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata13_w;
			end
			4'd9: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata12_w;
			end
			4'd10: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata11_w;
			end
			4'd11: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata10_w;
			end
			4'd12: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata9_w;
			end
			4'd13: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata8_w;
			end
			4'd14: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata7_w;
			end
			4'd15: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata6_w;
			end
			5'd16: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata5_w;
			end
			5'd17: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata4_w;
			end
			5'd18: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata3_w;
			end
			5'd19: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata2_w;
			end
			5'd20: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata1_w;
			end
			5'd21: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_wrdata0_w;
			end
			5'd22: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata15_w;
			end
			5'd23: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata14_w;
			end
			5'd24: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata13_w;
			end
			5'd25: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata12_w;
			end
			5'd26: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata11_w;
			end
			5'd27: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata10_w;
			end
			5'd28: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata9_w;
			end
			5'd29: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata8_w;
			end
			5'd30: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata7_w;
			end
			5'd31: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata6_w;
			end
			6'd32: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata5_w;
			end
			6'd33: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata4_w;
			end
			6'd34: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata3_w;
			end
			6'd35: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata2_w;
			end
			6'd36: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata1_w;
			end
			6'd37: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi0_rddata0_w;
			end
			6'd38: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_command0_w;
			end
			6'd39: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= main_nist_clock_nist_clock_phaseinjector1_command_issue_w;
			end
			6'd40: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_address1_w;
			end
			6'd41: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_address0_w;
			end
			6'd42: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_baddress0_w;
			end
			6'd43: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata15_w;
			end
			6'd44: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata14_w;
			end
			6'd45: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata13_w;
			end
			6'd46: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata12_w;
			end
			6'd47: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata11_w;
			end
			6'd48: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata10_w;
			end
			6'd49: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata9_w;
			end
			6'd50: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata8_w;
			end
			6'd51: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata7_w;
			end
			6'd52: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata6_w;
			end
			6'd53: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata5_w;
			end
			6'd54: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata4_w;
			end
			6'd55: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata3_w;
			end
			6'd56: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata2_w;
			end
			6'd57: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata1_w;
			end
			6'd58: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_wrdata0_w;
			end
			6'd59: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata15_w;
			end
			6'd60: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata14_w;
			end
			6'd61: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata13_w;
			end
			6'd62: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata12_w;
			end
			6'd63: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata11_w;
			end
			7'd64: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata10_w;
			end
			7'd65: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata9_w;
			end
			7'd66: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata8_w;
			end
			7'd67: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata7_w;
			end
			7'd68: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata6_w;
			end
			7'd69: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata5_w;
			end
			7'd70: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata4_w;
			end
			7'd71: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata3_w;
			end
			7'd72: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata2_w;
			end
			7'd73: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata1_w;
			end
			7'd74: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi1_rddata0_w;
			end
			7'd75: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_command0_w;
			end
			7'd76: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= main_nist_clock_nist_clock_phaseinjector2_command_issue_w;
			end
			7'd77: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_address1_w;
			end
			7'd78: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_address0_w;
			end
			7'd79: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_baddress0_w;
			end
			7'd80: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata15_w;
			end
			7'd81: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata14_w;
			end
			7'd82: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata13_w;
			end
			7'd83: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata12_w;
			end
			7'd84: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata11_w;
			end
			7'd85: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata10_w;
			end
			7'd86: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata9_w;
			end
			7'd87: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata8_w;
			end
			7'd88: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata7_w;
			end
			7'd89: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata6_w;
			end
			7'd90: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata5_w;
			end
			7'd91: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata4_w;
			end
			7'd92: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata3_w;
			end
			7'd93: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata2_w;
			end
			7'd94: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata1_w;
			end
			7'd95: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_wrdata0_w;
			end
			7'd96: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata15_w;
			end
			7'd97: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata14_w;
			end
			7'd98: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata13_w;
			end
			7'd99: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata12_w;
			end
			7'd100: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata11_w;
			end
			7'd101: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata10_w;
			end
			7'd102: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata9_w;
			end
			7'd103: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata8_w;
			end
			7'd104: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata7_w;
			end
			7'd105: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata6_w;
			end
			7'd106: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata5_w;
			end
			7'd107: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata4_w;
			end
			7'd108: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata3_w;
			end
			7'd109: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata2_w;
			end
			7'd110: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata1_w;
			end
			7'd111: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi2_rddata0_w;
			end
			7'd112: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_command0_w;
			end
			7'd113: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= main_nist_clock_nist_clock_phaseinjector3_command_issue_w;
			end
			7'd114: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_address1_w;
			end
			7'd115: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_address0_w;
			end
			7'd116: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_baddress0_w;
			end
			7'd117: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata15_w;
			end
			7'd118: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata14_w;
			end
			7'd119: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata13_w;
			end
			7'd120: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata12_w;
			end
			7'd121: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata11_w;
			end
			7'd122: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata10_w;
			end
			7'd123: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata9_w;
			end
			7'd124: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata8_w;
			end
			7'd125: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata7_w;
			end
			7'd126: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata6_w;
			end
			7'd127: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata5_w;
			end
			8'd128: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata4_w;
			end
			8'd129: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata3_w;
			end
			8'd130: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata2_w;
			end
			8'd131: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata1_w;
			end
			8'd132: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_wrdata0_w;
			end
			8'd133: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata15_w;
			end
			8'd134: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata14_w;
			end
			8'd135: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata13_w;
			end
			8'd136: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata12_w;
			end
			8'd137: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata11_w;
			end
			8'd138: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata10_w;
			end
			8'd139: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata9_w;
			end
			8'd140: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata8_w;
			end
			8'd141: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata7_w;
			end
			8'd142: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata6_w;
			end
			8'd143: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata5_w;
			end
			8'd144: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata4_w;
			end
			8'd145: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata3_w;
			end
			8'd146: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata2_w;
			end
			8'd147: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata1_w;
			end
			8'd148: begin
				builder_nist_clock_interface1_bank_bus_dat_r <= builder_nist_clock_csrbank1_pi3_rddata0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank1_control0_re) begin
		main_nist_clock_nist_clock_storage_full[3:0] <= builder_nist_clock_csrbank1_control0_r;
	end
	main_nist_clock_nist_clock_re <= builder_nist_clock_csrbank1_control0_re;
	if (builder_nist_clock_csrbank1_pi0_command0_re) begin
		main_nist_clock_nist_clock_phaseinjector0_command_storage_full[5:0] <= builder_nist_clock_csrbank1_pi0_command0_r;
	end
	main_nist_clock_nist_clock_phaseinjector0_command_re <= builder_nist_clock_csrbank1_pi0_command0_re;
	if (builder_nist_clock_csrbank1_pi0_address1_re) begin
		main_nist_clock_nist_clock_phaseinjector0_address_storage_full[13:8] <= builder_nist_clock_csrbank1_pi0_address1_r;
	end
	if (builder_nist_clock_csrbank1_pi0_address0_re) begin
		main_nist_clock_nist_clock_phaseinjector0_address_storage_full[7:0] <= builder_nist_clock_csrbank1_pi0_address0_r;
	end
	main_nist_clock_nist_clock_phaseinjector0_address_re <= builder_nist_clock_csrbank1_pi0_address0_re;
	if (builder_nist_clock_csrbank1_pi0_baddress0_re) begin
		main_nist_clock_nist_clock_phaseinjector0_baddress_storage_full[2:0] <= builder_nist_clock_csrbank1_pi0_baddress0_r;
	end
	main_nist_clock_nist_clock_phaseinjector0_baddress_re <= builder_nist_clock_csrbank1_pi0_baddress0_re;
	if (builder_nist_clock_csrbank1_pi0_wrdata15_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[127:120] <= builder_nist_clock_csrbank1_pi0_wrdata15_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata14_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[119:112] <= builder_nist_clock_csrbank1_pi0_wrdata14_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata13_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[111:104] <= builder_nist_clock_csrbank1_pi0_wrdata13_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata12_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[103:96] <= builder_nist_clock_csrbank1_pi0_wrdata12_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata11_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[95:88] <= builder_nist_clock_csrbank1_pi0_wrdata11_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata10_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[87:80] <= builder_nist_clock_csrbank1_pi0_wrdata10_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata9_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[79:72] <= builder_nist_clock_csrbank1_pi0_wrdata9_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata8_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[71:64] <= builder_nist_clock_csrbank1_pi0_wrdata8_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata7_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[63:56] <= builder_nist_clock_csrbank1_pi0_wrdata7_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata6_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[55:48] <= builder_nist_clock_csrbank1_pi0_wrdata6_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata5_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[47:40] <= builder_nist_clock_csrbank1_pi0_wrdata5_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata4_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[39:32] <= builder_nist_clock_csrbank1_pi0_wrdata4_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata3_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[31:24] <= builder_nist_clock_csrbank1_pi0_wrdata3_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata2_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[23:16] <= builder_nist_clock_csrbank1_pi0_wrdata2_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata1_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[15:8] <= builder_nist_clock_csrbank1_pi0_wrdata1_r;
	end
	if (builder_nist_clock_csrbank1_pi0_wrdata0_re) begin
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full[7:0] <= builder_nist_clock_csrbank1_pi0_wrdata0_r;
	end
	main_nist_clock_nist_clock_phaseinjector0_wrdata_re <= builder_nist_clock_csrbank1_pi0_wrdata0_re;
	if (builder_nist_clock_csrbank1_pi1_command0_re) begin
		main_nist_clock_nist_clock_phaseinjector1_command_storage_full[5:0] <= builder_nist_clock_csrbank1_pi1_command0_r;
	end
	main_nist_clock_nist_clock_phaseinjector1_command_re <= builder_nist_clock_csrbank1_pi1_command0_re;
	if (builder_nist_clock_csrbank1_pi1_address1_re) begin
		main_nist_clock_nist_clock_phaseinjector1_address_storage_full[13:8] <= builder_nist_clock_csrbank1_pi1_address1_r;
	end
	if (builder_nist_clock_csrbank1_pi1_address0_re) begin
		main_nist_clock_nist_clock_phaseinjector1_address_storage_full[7:0] <= builder_nist_clock_csrbank1_pi1_address0_r;
	end
	main_nist_clock_nist_clock_phaseinjector1_address_re <= builder_nist_clock_csrbank1_pi1_address0_re;
	if (builder_nist_clock_csrbank1_pi1_baddress0_re) begin
		main_nist_clock_nist_clock_phaseinjector1_baddress_storage_full[2:0] <= builder_nist_clock_csrbank1_pi1_baddress0_r;
	end
	main_nist_clock_nist_clock_phaseinjector1_baddress_re <= builder_nist_clock_csrbank1_pi1_baddress0_re;
	if (builder_nist_clock_csrbank1_pi1_wrdata15_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[127:120] <= builder_nist_clock_csrbank1_pi1_wrdata15_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata14_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[119:112] <= builder_nist_clock_csrbank1_pi1_wrdata14_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata13_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[111:104] <= builder_nist_clock_csrbank1_pi1_wrdata13_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata12_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[103:96] <= builder_nist_clock_csrbank1_pi1_wrdata12_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata11_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[95:88] <= builder_nist_clock_csrbank1_pi1_wrdata11_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata10_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[87:80] <= builder_nist_clock_csrbank1_pi1_wrdata10_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata9_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[79:72] <= builder_nist_clock_csrbank1_pi1_wrdata9_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata8_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[71:64] <= builder_nist_clock_csrbank1_pi1_wrdata8_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata7_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[63:56] <= builder_nist_clock_csrbank1_pi1_wrdata7_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata6_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[55:48] <= builder_nist_clock_csrbank1_pi1_wrdata6_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata5_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[47:40] <= builder_nist_clock_csrbank1_pi1_wrdata5_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata4_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[39:32] <= builder_nist_clock_csrbank1_pi1_wrdata4_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata3_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[31:24] <= builder_nist_clock_csrbank1_pi1_wrdata3_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata2_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[23:16] <= builder_nist_clock_csrbank1_pi1_wrdata2_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata1_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[15:8] <= builder_nist_clock_csrbank1_pi1_wrdata1_r;
	end
	if (builder_nist_clock_csrbank1_pi1_wrdata0_re) begin
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full[7:0] <= builder_nist_clock_csrbank1_pi1_wrdata0_r;
	end
	main_nist_clock_nist_clock_phaseinjector1_wrdata_re <= builder_nist_clock_csrbank1_pi1_wrdata0_re;
	if (builder_nist_clock_csrbank1_pi2_command0_re) begin
		main_nist_clock_nist_clock_phaseinjector2_command_storage_full[5:0] <= builder_nist_clock_csrbank1_pi2_command0_r;
	end
	main_nist_clock_nist_clock_phaseinjector2_command_re <= builder_nist_clock_csrbank1_pi2_command0_re;
	if (builder_nist_clock_csrbank1_pi2_address1_re) begin
		main_nist_clock_nist_clock_phaseinjector2_address_storage_full[13:8] <= builder_nist_clock_csrbank1_pi2_address1_r;
	end
	if (builder_nist_clock_csrbank1_pi2_address0_re) begin
		main_nist_clock_nist_clock_phaseinjector2_address_storage_full[7:0] <= builder_nist_clock_csrbank1_pi2_address0_r;
	end
	main_nist_clock_nist_clock_phaseinjector2_address_re <= builder_nist_clock_csrbank1_pi2_address0_re;
	if (builder_nist_clock_csrbank1_pi2_baddress0_re) begin
		main_nist_clock_nist_clock_phaseinjector2_baddress_storage_full[2:0] <= builder_nist_clock_csrbank1_pi2_baddress0_r;
	end
	main_nist_clock_nist_clock_phaseinjector2_baddress_re <= builder_nist_clock_csrbank1_pi2_baddress0_re;
	if (builder_nist_clock_csrbank1_pi2_wrdata15_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[127:120] <= builder_nist_clock_csrbank1_pi2_wrdata15_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata14_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[119:112] <= builder_nist_clock_csrbank1_pi2_wrdata14_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata13_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[111:104] <= builder_nist_clock_csrbank1_pi2_wrdata13_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata12_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[103:96] <= builder_nist_clock_csrbank1_pi2_wrdata12_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata11_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[95:88] <= builder_nist_clock_csrbank1_pi2_wrdata11_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata10_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[87:80] <= builder_nist_clock_csrbank1_pi2_wrdata10_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata9_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[79:72] <= builder_nist_clock_csrbank1_pi2_wrdata9_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata8_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[71:64] <= builder_nist_clock_csrbank1_pi2_wrdata8_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata7_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[63:56] <= builder_nist_clock_csrbank1_pi2_wrdata7_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata6_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[55:48] <= builder_nist_clock_csrbank1_pi2_wrdata6_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata5_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[47:40] <= builder_nist_clock_csrbank1_pi2_wrdata5_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata4_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[39:32] <= builder_nist_clock_csrbank1_pi2_wrdata4_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata3_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[31:24] <= builder_nist_clock_csrbank1_pi2_wrdata3_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata2_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[23:16] <= builder_nist_clock_csrbank1_pi2_wrdata2_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata1_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[15:8] <= builder_nist_clock_csrbank1_pi2_wrdata1_r;
	end
	if (builder_nist_clock_csrbank1_pi2_wrdata0_re) begin
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full[7:0] <= builder_nist_clock_csrbank1_pi2_wrdata0_r;
	end
	main_nist_clock_nist_clock_phaseinjector2_wrdata_re <= builder_nist_clock_csrbank1_pi2_wrdata0_re;
	if (builder_nist_clock_csrbank1_pi3_command0_re) begin
		main_nist_clock_nist_clock_phaseinjector3_command_storage_full[5:0] <= builder_nist_clock_csrbank1_pi3_command0_r;
	end
	main_nist_clock_nist_clock_phaseinjector3_command_re <= builder_nist_clock_csrbank1_pi3_command0_re;
	if (builder_nist_clock_csrbank1_pi3_address1_re) begin
		main_nist_clock_nist_clock_phaseinjector3_address_storage_full[13:8] <= builder_nist_clock_csrbank1_pi3_address1_r;
	end
	if (builder_nist_clock_csrbank1_pi3_address0_re) begin
		main_nist_clock_nist_clock_phaseinjector3_address_storage_full[7:0] <= builder_nist_clock_csrbank1_pi3_address0_r;
	end
	main_nist_clock_nist_clock_phaseinjector3_address_re <= builder_nist_clock_csrbank1_pi3_address0_re;
	if (builder_nist_clock_csrbank1_pi3_baddress0_re) begin
		main_nist_clock_nist_clock_phaseinjector3_baddress_storage_full[2:0] <= builder_nist_clock_csrbank1_pi3_baddress0_r;
	end
	main_nist_clock_nist_clock_phaseinjector3_baddress_re <= builder_nist_clock_csrbank1_pi3_baddress0_re;
	if (builder_nist_clock_csrbank1_pi3_wrdata15_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[127:120] <= builder_nist_clock_csrbank1_pi3_wrdata15_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata14_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[119:112] <= builder_nist_clock_csrbank1_pi3_wrdata14_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata13_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[111:104] <= builder_nist_clock_csrbank1_pi3_wrdata13_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata12_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[103:96] <= builder_nist_clock_csrbank1_pi3_wrdata12_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata11_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[95:88] <= builder_nist_clock_csrbank1_pi3_wrdata11_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata10_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[87:80] <= builder_nist_clock_csrbank1_pi3_wrdata10_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata9_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[79:72] <= builder_nist_clock_csrbank1_pi3_wrdata9_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata8_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[71:64] <= builder_nist_clock_csrbank1_pi3_wrdata8_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata7_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[63:56] <= builder_nist_clock_csrbank1_pi3_wrdata7_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata6_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[55:48] <= builder_nist_clock_csrbank1_pi3_wrdata6_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata5_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[47:40] <= builder_nist_clock_csrbank1_pi3_wrdata5_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata4_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[39:32] <= builder_nist_clock_csrbank1_pi3_wrdata4_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata3_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[31:24] <= builder_nist_clock_csrbank1_pi3_wrdata3_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata2_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[23:16] <= builder_nist_clock_csrbank1_pi3_wrdata2_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata1_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[15:8] <= builder_nist_clock_csrbank1_pi3_wrdata1_r;
	end
	if (builder_nist_clock_csrbank1_pi3_wrdata0_re) begin
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full[7:0] <= builder_nist_clock_csrbank1_pi3_wrdata0_r;
	end
	main_nist_clock_nist_clock_phaseinjector3_wrdata_re <= builder_nist_clock_csrbank1_pi3_wrdata0_re;
	builder_nist_clock_interface2_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank2_sel) begin
		case (builder_nist_clock_interface2_bank_bus_adr[4:0])
			1'd0: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_slot_w;
			end
			1'd1: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_length3_w;
			end
			2'd2: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_length2_w;
			end
			2'd3: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_length1_w;
			end
			3'd4: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_length0_w;
			end
			3'd5: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_errors3_w;
			end
			3'd6: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_errors2_w;
			end
			3'd7: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_errors1_w;
			end
			4'd8: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_errors0_w;
			end
			4'd9: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= main_writer_status_w;
			end
			4'd10: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= main_writer_pending_w;
			end
			4'd11: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_writer_ev_enable0_w;
			end
			4'd12: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= main_reader_start_w;
			end
			4'd13: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_reader_ready_w;
			end
			4'd14: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_reader_slot0_w;
			end
			4'd15: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_reader_length1_w;
			end
			5'd16: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_reader_length0_w;
			end
			5'd17: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= main_reader_eventmanager_status_w;
			end
			5'd18: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= main_reader_eventmanager_pending_w;
			end
			5'd19: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_sram_reader_ev_enable0_w;
			end
			5'd20: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_preamble_errors3_w;
			end
			5'd21: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_preamble_errors2_w;
			end
			5'd22: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_preamble_errors1_w;
			end
			5'd23: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_preamble_errors0_w;
			end
			5'd24: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_crc_errors3_w;
			end
			5'd25: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_crc_errors2_w;
			end
			5'd26: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_crc_errors1_w;
			end
			5'd27: begin
				builder_nist_clock_interface2_bank_bus_dat_r <= builder_nist_clock_csrbank2_crc_errors0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank2_sram_writer_ev_enable0_re) begin
		main_writer_storage_full <= builder_nist_clock_csrbank2_sram_writer_ev_enable0_r;
	end
	main_writer_re <= builder_nist_clock_csrbank2_sram_writer_ev_enable0_re;
	if (builder_nist_clock_csrbank2_sram_reader_slot0_re) begin
		main_reader_slot_storage_full[1:0] <= builder_nist_clock_csrbank2_sram_reader_slot0_r;
	end
	main_reader_slot_re <= builder_nist_clock_csrbank2_sram_reader_slot0_re;
	if (builder_nist_clock_csrbank2_sram_reader_length1_re) begin
		main_reader_length_storage_full[10:8] <= builder_nist_clock_csrbank2_sram_reader_length1_r;
	end
	if (builder_nist_clock_csrbank2_sram_reader_length0_re) begin
		main_reader_length_storage_full[7:0] <= builder_nist_clock_csrbank2_sram_reader_length0_r;
	end
	main_reader_length_re <= builder_nist_clock_csrbank2_sram_reader_length0_re;
	if (builder_nist_clock_csrbank2_sram_reader_ev_enable0_re) begin
		main_reader_eventmanager_storage_full <= builder_nist_clock_csrbank2_sram_reader_ev_enable0_r;
	end
	main_reader_eventmanager_re <= builder_nist_clock_csrbank2_sram_reader_ev_enable0_re;
	builder_nist_clock_interface3_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank3_sel) begin
		case (builder_nist_clock_interface3_bank_bus_adr[0])
			1'd0: begin
				builder_nist_clock_interface3_bank_bus_dat_r <= builder_nist_clock_csrbank3_mode_detection_mode_w;
			end
			1'd1: begin
				builder_nist_clock_interface3_bank_bus_dat_r <= builder_nist_clock_csrbank3_crg_reset0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank3_crg_reset0_re) begin
		main_ethphy_storage_full <= builder_nist_clock_csrbank3_crg_reset0_r;
	end
	main_ethphy_re <= builder_nist_clock_csrbank3_crg_reset0_re;
	builder_nist_clock_interface4_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank4_sel) begin
		case (builder_nist_clock_interface4_bank_bus_adr[1:0])
			1'd0: begin
				builder_nist_clock_interface4_bank_bus_dat_r <= builder_nist_clock_csrbank4_in_w;
			end
			1'd1: begin
				builder_nist_clock_interface4_bank_bus_dat_r <= builder_nist_clock_csrbank4_out0_w;
			end
			2'd2: begin
				builder_nist_clock_interface4_bank_bus_dat_r <= builder_nist_clock_csrbank4_oe0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank4_out0_re) begin
		main_i2c_out_storage_full[1:0] <= builder_nist_clock_csrbank4_out0_r;
	end
	main_i2c_out_re <= builder_nist_clock_csrbank4_out0_re;
	if (builder_nist_clock_csrbank4_oe0_re) begin
		main_i2c_oe_storage_full[1:0] <= builder_nist_clock_csrbank4_oe0_r;
	end
	main_i2c_oe_re <= builder_nist_clock_csrbank4_oe0_re;
	builder_nist_clock_interface5_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank5_sel) begin
		case (builder_nist_clock_interface5_bank_bus_adr[0])
			1'd0: begin
				builder_nist_clock_interface5_bank_bus_dat_r <= builder_nist_clock_csrbank5_address0_w;
			end
			1'd1: begin
				builder_nist_clock_interface5_bank_bus_dat_r <= builder_nist_clock_csrbank5_data_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank5_address0_re) begin
		main_add_identifier_storage_full[7:0] <= builder_nist_clock_csrbank5_address0_r;
	end
	main_add_identifier_re <= builder_nist_clock_csrbank5_address0_re;
	builder_nist_clock_interface6_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank6_sel) begin
		case (builder_nist_clock_interface6_bank_bus_adr[0])
			1'd0: begin
				builder_nist_clock_interface6_bank_bus_dat_r <= builder_nist_clock_csrbank6_reset0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank6_reset0_re) begin
		main_kernel_cpu_storage_full <= builder_nist_clock_csrbank6_reset0_r;
	end
	main_kernel_cpu_re <= builder_nist_clock_csrbank6_reset0_re;
	builder_nist_clock_interface7_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank7_sel) begin
		case (builder_nist_clock_interface7_bank_bus_adr[0])
			1'd0: begin
				builder_nist_clock_interface7_bank_bus_dat_r <= builder_nist_clock_csrbank7_out0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank7_out0_re) begin
		main_leds_storage_full[1:0] <= builder_nist_clock_csrbank7_out0_r;
	end
	main_leds_re <= builder_nist_clock_csrbank7_out0_re;
	builder_nist_clock_interface8_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank8_sel) begin
		case (builder_nist_clock_interface8_bank_bus_adr[4:0])
			1'd0: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_enable0_w;
			end
			1'd1: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_busy_w;
			end
			2'd2: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_message_encoder_overflow_w;
			end
			2'd3: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= main_rtio_analyzer_message_encoder_overflow_reset_w;
			end
			3'd4: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= main_rtio_analyzer_dma_reset_w;
			end
			3'd5: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_base_address4_w;
			end
			3'd6: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_base_address3_w;
			end
			3'd7: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_base_address2_w;
			end
			4'd8: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_base_address1_w;
			end
			4'd9: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_base_address0_w;
			end
			4'd10: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_last_address4_w;
			end
			4'd11: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_last_address3_w;
			end
			4'd12: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_last_address2_w;
			end
			4'd13: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_last_address1_w;
			end
			4'd14: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_last_address0_w;
			end
			4'd15: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count7_w;
			end
			5'd16: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count6_w;
			end
			5'd17: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count5_w;
			end
			5'd18: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count4_w;
			end
			5'd19: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count3_w;
			end
			5'd20: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count2_w;
			end
			5'd21: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count1_w;
			end
			5'd22: begin
				builder_nist_clock_interface8_bank_bus_dat_r <= builder_nist_clock_csrbank8_dma_byte_count0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank8_enable0_re) begin
		main_rtio_analyzer_enable_storage_full <= builder_nist_clock_csrbank8_enable0_r;
	end
	main_rtio_analyzer_enable_re <= builder_nist_clock_csrbank8_enable0_re;
	if (builder_nist_clock_csrbank8_dma_base_address4_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[35:32] <= builder_nist_clock_csrbank8_dma_base_address4_r;
	end
	if (builder_nist_clock_csrbank8_dma_base_address3_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[31:24] <= builder_nist_clock_csrbank8_dma_base_address3_r;
	end
	if (builder_nist_clock_csrbank8_dma_base_address2_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[23:16] <= builder_nist_clock_csrbank8_dma_base_address2_r;
	end
	if (builder_nist_clock_csrbank8_dma_base_address1_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[15:8] <= builder_nist_clock_csrbank8_dma_base_address1_r;
	end
	if (builder_nist_clock_csrbank8_dma_base_address0_re) begin
		main_rtio_analyzer_dma_base_address_storage_full[7:0] <= builder_nist_clock_csrbank8_dma_base_address0_r;
	end
	main_rtio_analyzer_dma_base_address_re <= builder_nist_clock_csrbank8_dma_base_address0_re;
	if (builder_nist_clock_csrbank8_dma_last_address4_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[35:32] <= builder_nist_clock_csrbank8_dma_last_address4_r;
	end
	if (builder_nist_clock_csrbank8_dma_last_address3_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[31:24] <= builder_nist_clock_csrbank8_dma_last_address3_r;
	end
	if (builder_nist_clock_csrbank8_dma_last_address2_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[23:16] <= builder_nist_clock_csrbank8_dma_last_address2_r;
	end
	if (builder_nist_clock_csrbank8_dma_last_address1_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[15:8] <= builder_nist_clock_csrbank8_dma_last_address1_r;
	end
	if (builder_nist_clock_csrbank8_dma_last_address0_re) begin
		main_rtio_analyzer_dma_last_address_storage_full[7:0] <= builder_nist_clock_csrbank8_dma_last_address0_r;
	end
	main_rtio_analyzer_dma_last_address_re <= builder_nist_clock_csrbank8_dma_last_address0_re;
	builder_nist_clock_interface9_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank9_sel) begin
		case (builder_nist_clock_interface9_bank_bus_adr[3:0])
			1'd0: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= main_rtio_core_reset_w;
			end
			1'd1: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= main_rtio_core_reset_phy_w;
			end
			2'd2: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= main_rtio_core_async_error_w;
			end
			2'd3: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_collision_channel1_w;
			end
			3'd4: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_collision_channel0_w;
			end
			3'd5: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_busy_channel1_w;
			end
			3'd6: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_busy_channel0_w;
			end
			3'd7: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_sequence_error_channel1_w;
			end
			4'd8: begin
				builder_nist_clock_interface9_bank_bus_dat_r <= builder_nist_clock_csrbank9_sequence_error_channel0_w;
			end
		endcase
	end
	builder_nist_clock_interface10_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank10_sel) begin
		case (builder_nist_clock_interface10_bank_bus_adr[1:0])
			1'd0: begin
				builder_nist_clock_interface10_bank_bus_dat_r <= builder_nist_clock_csrbank10_clock_sel0_w;
			end
			1'd1: begin
				builder_nist_clock_interface10_bank_bus_dat_r <= builder_nist_clock_csrbank10_pll_reset0_w;
			end
			2'd2: begin
				builder_nist_clock_interface10_bank_bus_dat_r <= builder_nist_clock_csrbank10_pll_locked_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank10_clock_sel0_re) begin
		main_rtio_crg_clock_sel_storage_full <= builder_nist_clock_csrbank10_clock_sel0_r;
	end
	main_rtio_crg_clock_sel_re <= builder_nist_clock_csrbank10_clock_sel0_re;
	if (builder_nist_clock_csrbank10_pll_reset0_re) begin
		main_rtio_crg_pll_reset_storage_full <= builder_nist_clock_csrbank10_pll_reset0_r;
	end
	main_rtio_crg_pll_reset_re <= builder_nist_clock_csrbank10_pll_reset0_re;
	builder_nist_clock_interface11_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank11_sel) begin
		case (builder_nist_clock_interface11_bank_bus_adr[3:0])
			1'd0: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_chan_sel0_w;
			end
			1'd1: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_probe_sel0_w;
			end
			2'd2: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= main_mon_value_update_w;
			end
			2'd3: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_value3_w;
			end
			3'd4: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_value2_w;
			end
			3'd5: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_value1_w;
			end
			3'd6: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_mon_value0_w;
			end
			3'd7: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_inj_chan_sel0_w;
			end
			4'd8: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= builder_nist_clock_csrbank11_inj_override_sel0_w;
			end
			4'd9: begin
				builder_nist_clock_interface11_bank_bus_dat_r <= main_inj_value_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank11_mon_chan_sel0_re) begin
		main_mon_chan_sel_storage_full[4:0] <= builder_nist_clock_csrbank11_mon_chan_sel0_r;
	end
	main_mon_chan_sel_re <= builder_nist_clock_csrbank11_mon_chan_sel0_re;
	if (builder_nist_clock_csrbank11_mon_probe_sel0_re) begin
		main_mon_probe_sel_storage_full[3:0] <= builder_nist_clock_csrbank11_mon_probe_sel0_r;
	end
	main_mon_probe_sel_re <= builder_nist_clock_csrbank11_mon_probe_sel0_re;
	if (builder_nist_clock_csrbank11_inj_chan_sel0_re) begin
		main_inj_chan_sel_storage_full[4:0] <= builder_nist_clock_csrbank11_inj_chan_sel0_r;
	end
	main_inj_chan_sel_re <= builder_nist_clock_csrbank11_inj_chan_sel0_re;
	if (builder_nist_clock_csrbank11_inj_override_sel0_re) begin
		main_inj_override_sel_storage_full[1:0] <= builder_nist_clock_csrbank11_inj_override_sel0_r;
	end
	main_inj_override_sel_re <= builder_nist_clock_csrbank11_inj_override_sel0_re;
	builder_nist_clock_interface12_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank12_sel) begin
		case (builder_nist_clock_interface12_bank_bus_adr[1:0])
			1'd0: begin
				builder_nist_clock_interface12_bank_bus_dat_r <= builder_nist_clock_csrbank12_bitbang0_w;
			end
			1'd1: begin
				builder_nist_clock_interface12_bank_bus_dat_r <= builder_nist_clock_csrbank12_miso_w;
			end
			2'd2: begin
				builder_nist_clock_interface12_bank_bus_dat_r <= builder_nist_clock_csrbank12_bitbang_en0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank12_bitbang0_re) begin
		main_nist_clock_spiflash_bitbang_storage_full[3:0] <= builder_nist_clock_csrbank12_bitbang0_r;
	end
	main_nist_clock_spiflash_bitbang_re <= builder_nist_clock_csrbank12_bitbang0_re;
	if (builder_nist_clock_csrbank12_bitbang_en0_re) begin
		main_nist_clock_spiflash_bitbang_en_storage_full <= builder_nist_clock_csrbank12_bitbang_en0_r;
	end
	main_nist_clock_spiflash_bitbang_en_re <= builder_nist_clock_csrbank12_bitbang_en0_re;
	builder_nist_clock_interface13_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank13_sel) begin
		case (builder_nist_clock_interface13_bank_bus_adr[4:0])
			1'd0: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load7_w;
			end
			1'd1: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load6_w;
			end
			2'd2: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load5_w;
			end
			2'd3: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load4_w;
			end
			3'd4: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load3_w;
			end
			3'd5: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load2_w;
			end
			3'd6: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load1_w;
			end
			3'd7: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_load0_w;
			end
			4'd8: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload7_w;
			end
			4'd9: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload6_w;
			end
			4'd10: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload5_w;
			end
			4'd11: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload4_w;
			end
			4'd12: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload3_w;
			end
			4'd13: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload2_w;
			end
			4'd14: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload1_w;
			end
			4'd15: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_reload0_w;
			end
			5'd16: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_en0_w;
			end
			5'd17: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= main_nist_clock_nist_clock_timer0_update_value_w;
			end
			5'd18: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value7_w;
			end
			5'd19: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value6_w;
			end
			5'd20: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value5_w;
			end
			5'd21: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value4_w;
			end
			5'd22: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value3_w;
			end
			5'd23: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value2_w;
			end
			5'd24: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value1_w;
			end
			5'd25: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_value0_w;
			end
			5'd26: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= main_nist_clock_nist_clock_timer0_eventmanager_status_w;
			end
			5'd27: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= main_nist_clock_nist_clock_timer0_eventmanager_pending_w;
			end
			5'd28: begin
				builder_nist_clock_interface13_bank_bus_dat_r <= builder_nist_clock_csrbank13_ev_enable0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank13_load7_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[63:56] <= builder_nist_clock_csrbank13_load7_r;
	end
	if (builder_nist_clock_csrbank13_load6_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[55:48] <= builder_nist_clock_csrbank13_load6_r;
	end
	if (builder_nist_clock_csrbank13_load5_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[47:40] <= builder_nist_clock_csrbank13_load5_r;
	end
	if (builder_nist_clock_csrbank13_load4_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[39:32] <= builder_nist_clock_csrbank13_load4_r;
	end
	if (builder_nist_clock_csrbank13_load3_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[31:24] <= builder_nist_clock_csrbank13_load3_r;
	end
	if (builder_nist_clock_csrbank13_load2_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[23:16] <= builder_nist_clock_csrbank13_load2_r;
	end
	if (builder_nist_clock_csrbank13_load1_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[15:8] <= builder_nist_clock_csrbank13_load1_r;
	end
	if (builder_nist_clock_csrbank13_load0_re) begin
		main_nist_clock_nist_clock_timer0_load_storage_full[7:0] <= builder_nist_clock_csrbank13_load0_r;
	end
	main_nist_clock_nist_clock_timer0_load_re <= builder_nist_clock_csrbank13_load0_re;
	if (builder_nist_clock_csrbank13_reload7_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[63:56] <= builder_nist_clock_csrbank13_reload7_r;
	end
	if (builder_nist_clock_csrbank13_reload6_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[55:48] <= builder_nist_clock_csrbank13_reload6_r;
	end
	if (builder_nist_clock_csrbank13_reload5_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[47:40] <= builder_nist_clock_csrbank13_reload5_r;
	end
	if (builder_nist_clock_csrbank13_reload4_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[39:32] <= builder_nist_clock_csrbank13_reload4_r;
	end
	if (builder_nist_clock_csrbank13_reload3_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[31:24] <= builder_nist_clock_csrbank13_reload3_r;
	end
	if (builder_nist_clock_csrbank13_reload2_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[23:16] <= builder_nist_clock_csrbank13_reload2_r;
	end
	if (builder_nist_clock_csrbank13_reload1_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[15:8] <= builder_nist_clock_csrbank13_reload1_r;
	end
	if (builder_nist_clock_csrbank13_reload0_re) begin
		main_nist_clock_nist_clock_timer0_reload_storage_full[7:0] <= builder_nist_clock_csrbank13_reload0_r;
	end
	main_nist_clock_nist_clock_timer0_reload_re <= builder_nist_clock_csrbank13_reload0_re;
	if (builder_nist_clock_csrbank13_en0_re) begin
		main_nist_clock_nist_clock_timer0_en_storage_full <= builder_nist_clock_csrbank13_en0_r;
	end
	main_nist_clock_nist_clock_timer0_en_re <= builder_nist_clock_csrbank13_en0_re;
	if (builder_nist_clock_csrbank13_ev_enable0_re) begin
		main_nist_clock_nist_clock_timer0_eventmanager_storage_full <= builder_nist_clock_csrbank13_ev_enable0_r;
	end
	main_nist_clock_nist_clock_timer0_eventmanager_re <= builder_nist_clock_csrbank13_ev_enable0_re;
	builder_nist_clock_interface14_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank14_sel) begin
		case (builder_nist_clock_interface14_bank_bus_adr[4:0])
			1'd0: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load7_w;
			end
			1'd1: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load6_w;
			end
			2'd2: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load5_w;
			end
			2'd3: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load4_w;
			end
			3'd4: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load3_w;
			end
			3'd5: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load2_w;
			end
			3'd6: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load1_w;
			end
			3'd7: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_load0_w;
			end
			4'd8: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload7_w;
			end
			4'd9: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload6_w;
			end
			4'd10: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload5_w;
			end
			4'd11: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload4_w;
			end
			4'd12: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload3_w;
			end
			4'd13: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload2_w;
			end
			4'd14: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload1_w;
			end
			4'd15: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_reload0_w;
			end
			5'd16: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_en0_w;
			end
			5'd17: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= main_update_value_w;
			end
			5'd18: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value7_w;
			end
			5'd19: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value6_w;
			end
			5'd20: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value5_w;
			end
			5'd21: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value4_w;
			end
			5'd22: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value3_w;
			end
			5'd23: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value2_w;
			end
			5'd24: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value1_w;
			end
			5'd25: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_value0_w;
			end
			5'd26: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= main_eventmanager_status_w;
			end
			5'd27: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= main_eventmanager_pending_w;
			end
			5'd28: begin
				builder_nist_clock_interface14_bank_bus_dat_r <= builder_nist_clock_csrbank14_ev_enable0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank14_load7_re) begin
		main_load_storage_full[63:56] <= builder_nist_clock_csrbank14_load7_r;
	end
	if (builder_nist_clock_csrbank14_load6_re) begin
		main_load_storage_full[55:48] <= builder_nist_clock_csrbank14_load6_r;
	end
	if (builder_nist_clock_csrbank14_load5_re) begin
		main_load_storage_full[47:40] <= builder_nist_clock_csrbank14_load5_r;
	end
	if (builder_nist_clock_csrbank14_load4_re) begin
		main_load_storage_full[39:32] <= builder_nist_clock_csrbank14_load4_r;
	end
	if (builder_nist_clock_csrbank14_load3_re) begin
		main_load_storage_full[31:24] <= builder_nist_clock_csrbank14_load3_r;
	end
	if (builder_nist_clock_csrbank14_load2_re) begin
		main_load_storage_full[23:16] <= builder_nist_clock_csrbank14_load2_r;
	end
	if (builder_nist_clock_csrbank14_load1_re) begin
		main_load_storage_full[15:8] <= builder_nist_clock_csrbank14_load1_r;
	end
	if (builder_nist_clock_csrbank14_load0_re) begin
		main_load_storage_full[7:0] <= builder_nist_clock_csrbank14_load0_r;
	end
	main_load_re <= builder_nist_clock_csrbank14_load0_re;
	if (builder_nist_clock_csrbank14_reload7_re) begin
		main_reload_storage_full[63:56] <= builder_nist_clock_csrbank14_reload7_r;
	end
	if (builder_nist_clock_csrbank14_reload6_re) begin
		main_reload_storage_full[55:48] <= builder_nist_clock_csrbank14_reload6_r;
	end
	if (builder_nist_clock_csrbank14_reload5_re) begin
		main_reload_storage_full[47:40] <= builder_nist_clock_csrbank14_reload5_r;
	end
	if (builder_nist_clock_csrbank14_reload4_re) begin
		main_reload_storage_full[39:32] <= builder_nist_clock_csrbank14_reload4_r;
	end
	if (builder_nist_clock_csrbank14_reload3_re) begin
		main_reload_storage_full[31:24] <= builder_nist_clock_csrbank14_reload3_r;
	end
	if (builder_nist_clock_csrbank14_reload2_re) begin
		main_reload_storage_full[23:16] <= builder_nist_clock_csrbank14_reload2_r;
	end
	if (builder_nist_clock_csrbank14_reload1_re) begin
		main_reload_storage_full[15:8] <= builder_nist_clock_csrbank14_reload1_r;
	end
	if (builder_nist_clock_csrbank14_reload0_re) begin
		main_reload_storage_full[7:0] <= builder_nist_clock_csrbank14_reload0_r;
	end
	main_reload_re <= builder_nist_clock_csrbank14_reload0_re;
	if (builder_nist_clock_csrbank14_en0_re) begin
		main_en_storage_full <= builder_nist_clock_csrbank14_en0_r;
	end
	main_en_re <= builder_nist_clock_csrbank14_en0_re;
	if (builder_nist_clock_csrbank14_ev_enable0_re) begin
		main_eventmanager_storage_full <= builder_nist_clock_csrbank14_ev_enable0_r;
	end
	main_eventmanager_re <= builder_nist_clock_csrbank14_ev_enable0_re;
	builder_nist_clock_interface15_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank15_sel) begin
		case (builder_nist_clock_interface15_bank_bus_adr[2:0])
			1'd0: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_enable_null0_w;
			end
			1'd1: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_enable_prog0_w;
			end
			2'd2: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_prog_address3_w;
			end
			2'd3: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_prog_address2_w;
			end
			3'd4: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_prog_address1_w;
			end
			3'd5: begin
				builder_nist_clock_interface15_bank_bus_dat_r <= builder_nist_clock_csrbank15_prog_address0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank15_enable_null0_re) begin
		main_nist_clock_nist_clock_tmpu_enable_null_storage_full <= builder_nist_clock_csrbank15_enable_null0_r;
	end
	main_nist_clock_nist_clock_tmpu_enable_null_re <= builder_nist_clock_csrbank15_enable_null0_re;
	if (builder_nist_clock_csrbank15_enable_prog0_re) begin
		main_nist_clock_nist_clock_tmpu_enable_prog_storage_full <= builder_nist_clock_csrbank15_enable_prog0_r;
	end
	main_nist_clock_nist_clock_tmpu_enable_prog_re <= builder_nist_clock_csrbank15_enable_prog0_re;
	if (builder_nist_clock_csrbank15_prog_address3_re) begin
		main_nist_clock_nist_clock_tmpu_prog_address_storage_full[29:24] <= builder_nist_clock_csrbank15_prog_address3_r;
	end
	if (builder_nist_clock_csrbank15_prog_address2_re) begin
		main_nist_clock_nist_clock_tmpu_prog_address_storage_full[23:16] <= builder_nist_clock_csrbank15_prog_address2_r;
	end
	if (builder_nist_clock_csrbank15_prog_address1_re) begin
		main_nist_clock_nist_clock_tmpu_prog_address_storage_full[15:8] <= builder_nist_clock_csrbank15_prog_address1_r;
	end
	if (builder_nist_clock_csrbank15_prog_address0_re) begin
		main_nist_clock_nist_clock_tmpu_prog_address_storage_full[7:0] <= builder_nist_clock_csrbank15_prog_address0_r;
	end
	main_nist_clock_nist_clock_tmpu_prog_address_re <= builder_nist_clock_csrbank15_prog_address0_re;
	builder_nist_clock_interface16_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank16_sel) begin
		case (builder_nist_clock_interface16_bank_bus_adr[2:0])
			1'd0: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= main_nist_clock_nist_clock_uart_rxtx_w;
			end
			1'd1: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= builder_nist_clock_csrbank16_txfull_w;
			end
			2'd2: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= builder_nist_clock_csrbank16_rxempty_w;
			end
			2'd3: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= main_nist_clock_nist_clock_uart_status_w;
			end
			3'd4: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= main_nist_clock_nist_clock_uart_pending_w;
			end
			3'd5: begin
				builder_nist_clock_interface16_bank_bus_dat_r <= builder_nist_clock_csrbank16_ev_enable0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank16_ev_enable0_re) begin
		main_nist_clock_nist_clock_uart_storage_full[1:0] <= builder_nist_clock_csrbank16_ev_enable0_r;
	end
	main_nist_clock_nist_clock_uart_re <= builder_nist_clock_csrbank16_ev_enable0_re;
	builder_nist_clock_interface17_bank_bus_dat_r <= 1'd0;
	if (builder_nist_clock_csrbank17_sel) begin
		case (builder_nist_clock_interface17_bank_bus_adr[1:0])
			1'd0: begin
				builder_nist_clock_interface17_bank_bus_dat_r <= builder_nist_clock_csrbank17_tuning_word3_w;
			end
			1'd1: begin
				builder_nist_clock_interface17_bank_bus_dat_r <= builder_nist_clock_csrbank17_tuning_word2_w;
			end
			2'd2: begin
				builder_nist_clock_interface17_bank_bus_dat_r <= builder_nist_clock_csrbank17_tuning_word1_w;
			end
			2'd3: begin
				builder_nist_clock_interface17_bank_bus_dat_r <= builder_nist_clock_csrbank17_tuning_word0_w;
			end
		endcase
	end
	if (builder_nist_clock_csrbank17_tuning_word3_re) begin
		main_nist_clock_nist_clock_uart_phy_storage_full[31:24] <= builder_nist_clock_csrbank17_tuning_word3_r;
	end
	if (builder_nist_clock_csrbank17_tuning_word2_re) begin
		main_nist_clock_nist_clock_uart_phy_storage_full[23:16] <= builder_nist_clock_csrbank17_tuning_word2_r;
	end
	if (builder_nist_clock_csrbank17_tuning_word1_re) begin
		main_nist_clock_nist_clock_uart_phy_storage_full[15:8] <= builder_nist_clock_csrbank17_tuning_word1_r;
	end
	if (builder_nist_clock_csrbank17_tuning_word0_re) begin
		main_nist_clock_nist_clock_uart_phy_storage_full[7:0] <= builder_nist_clock_csrbank17_tuning_word0_r;
	end
	main_nist_clock_nist_clock_uart_phy_re <= builder_nist_clock_csrbank17_tuning_word0_re;
	if (sys_rst) begin
		main_nist_clock_nist_clock_tmpu_enable_null_storage_full <= 1'd0;
		main_nist_clock_nist_clock_tmpu_enable_null_re <= 1'd0;
		main_nist_clock_nist_clock_tmpu_enable_prog_storage_full <= 1'd0;
		main_nist_clock_nist_clock_tmpu_enable_prog_re <= 1'd0;
		main_nist_clock_nist_clock_tmpu_prog_address_storage_full <= 30'd0;
		main_nist_clock_nist_clock_tmpu_prog_address_re <= 1'd0;
		main_nist_clock_nist_clock_tmpu_error <= 1'd0;
		main_nist_clock_nist_clock_sram_bus_ack <= 1'd0;
		main_nist_clock_nist_clock_interface_adr <= 14'd0;
		main_nist_clock_nist_clock_interface_we <= 1'd0;
		main_nist_clock_nist_clock_interface_dat_w <= 8'd0;
		main_nist_clock_nist_clock_bus_wishbone_dat_r <= 32'd0;
		main_nist_clock_nist_clock_bus_wishbone_ack <= 1'd0;
		main_nist_clock_nist_clock_counter <= 2'd0;
		serial_tx <= 1'd1;
		main_nist_clock_nist_clock_uart_phy_storage_full <= 32'd3958241;
		main_nist_clock_nist_clock_uart_phy_re <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_sink_ack <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_uart_clk_txen <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_phase_accumulator_tx <= 32'd0;
		main_nist_clock_nist_clock_uart_phy_tx_reg <= 8'd0;
		main_nist_clock_nist_clock_uart_phy_tx_bitcount <= 4'd0;
		main_nist_clock_nist_clock_uart_phy_tx_busy <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_source_stb <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_source_payload_data <= 8'd0;
		main_nist_clock_nist_clock_uart_phy_uart_clk_rxen <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_phase_accumulator_rx <= 32'd0;
		main_nist_clock_nist_clock_uart_phy_rx_r <= 1'd0;
		main_nist_clock_nist_clock_uart_phy_rx_reg <= 8'd0;
		main_nist_clock_nist_clock_uart_phy_rx_bitcount <= 4'd0;
		main_nist_clock_nist_clock_uart_phy_rx_busy <= 1'd0;
		main_nist_clock_nist_clock_uart_tx_pending <= 1'd0;
		main_nist_clock_nist_clock_uart_tx_old_trigger <= 1'd0;
		main_nist_clock_nist_clock_uart_rx_pending <= 1'd0;
		main_nist_clock_nist_clock_uart_rx_old_trigger <= 1'd0;
		main_nist_clock_nist_clock_uart_storage_full <= 2'd0;
		main_nist_clock_nist_clock_uart_re <= 1'd0;
		main_nist_clock_nist_clock_uart_tx_fifo_level <= 5'd0;
		main_nist_clock_nist_clock_uart_tx_fifo_produce <= 4'd0;
		main_nist_clock_nist_clock_uart_tx_fifo_consume <= 4'd0;
		main_nist_clock_nist_clock_uart_rx_fifo_level <= 5'd0;
		main_nist_clock_nist_clock_uart_rx_fifo_produce <= 4'd0;
		main_nist_clock_nist_clock_uart_rx_fifo_consume <= 4'd0;
		main_nist_clock_nist_clock_timer0_load_storage_full <= 64'd0;
		main_nist_clock_nist_clock_timer0_load_re <= 1'd0;
		main_nist_clock_nist_clock_timer0_reload_storage_full <= 64'd0;
		main_nist_clock_nist_clock_timer0_reload_re <= 1'd0;
		main_nist_clock_nist_clock_timer0_en_storage_full <= 1'd0;
		main_nist_clock_nist_clock_timer0_en_re <= 1'd0;
		main_nist_clock_nist_clock_timer0_value_status <= 64'd0;
		main_nist_clock_nist_clock_timer0_zero_pending <= 1'd0;
		main_nist_clock_nist_clock_timer0_zero_old_trigger <= 1'd0;
		main_nist_clock_nist_clock_timer0_eventmanager_storage_full <= 1'd0;
		main_nist_clock_nist_clock_timer0_eventmanager_re <= 1'd0;
		main_nist_clock_nist_clock_timer0_value <= 64'd0;
		main_nist_clock_ddrphy_wlevel_en_storage_full <= 1'd0;
		main_nist_clock_ddrphy_wlevel_en_re <= 1'd0;
		main_nist_clock_ddrphy_dly_sel_storage_full <= 8'd0;
		main_nist_clock_ddrphy_dly_sel_re <= 1'd0;
		main_nist_clock_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		main_nist_clock_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		main_nist_clock_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		main_nist_clock_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		main_nist_clock_ddrphy_oe_dqs <= 1'd0;
		main_nist_clock_ddrphy_oe_dq <= 1'd0;
		main_nist_clock_ddrphy_n_rddata_en0 <= 1'd0;
		main_nist_clock_ddrphy_n_rddata_en1 <= 1'd0;
		main_nist_clock_ddrphy_n_rddata_en2 <= 1'd0;
		main_nist_clock_ddrphy_n_rddata_en3 <= 1'd0;
		main_nist_clock_ddrphy_n_rddata_en4 <= 1'd0;
		main_nist_clock_ddrphy_last_wrdata_en <= 4'd0;
		main_nist_clock_nist_clock_storage_full <= 4'd0;
		main_nist_clock_nist_clock_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector0_command_storage_full <= 6'd0;
		main_nist_clock_nist_clock_phaseinjector0_command_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector0_address_storage_full <= 14'd0;
		main_nist_clock_nist_clock_phaseinjector0_address_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector0_baddress_storage_full <= 3'd0;
		main_nist_clock_nist_clock_phaseinjector0_baddress_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector0_wrdata_storage_full <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector0_wrdata_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector0_status <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector1_command_storage_full <= 6'd0;
		main_nist_clock_nist_clock_phaseinjector1_command_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector1_address_storage_full <= 14'd0;
		main_nist_clock_nist_clock_phaseinjector1_address_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector1_baddress_storage_full <= 3'd0;
		main_nist_clock_nist_clock_phaseinjector1_baddress_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector1_wrdata_storage_full <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector1_wrdata_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector1_status <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector2_command_storage_full <= 6'd0;
		main_nist_clock_nist_clock_phaseinjector2_command_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector2_address_storage_full <= 14'd0;
		main_nist_clock_nist_clock_phaseinjector2_address_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector2_baddress_storage_full <= 3'd0;
		main_nist_clock_nist_clock_phaseinjector2_baddress_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector2_wrdata_storage_full <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector2_wrdata_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector2_status <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector3_command_storage_full <= 6'd0;
		main_nist_clock_nist_clock_phaseinjector3_command_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector3_address_storage_full <= 14'd0;
		main_nist_clock_nist_clock_phaseinjector3_address_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector3_baddress_storage_full <= 3'd0;
		main_nist_clock_nist_clock_phaseinjector3_baddress_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector3_wrdata_storage_full <= 128'd0;
		main_nist_clock_nist_clock_phaseinjector3_wrdata_re <= 1'd0;
		main_nist_clock_nist_clock_phaseinjector3_status <= 128'd0;
		main_nist_clock_nist_clock_sdram_controller_bank0_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank0_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank1_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank1_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank2_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank2_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank3_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank3_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank4_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank4_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank5_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank5_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank6_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank6_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_bank7_idle <= 1'd1;
		main_nist_clock_nist_clock_sdram_controller_bank7_row1 <= 14'd0;
		main_nist_clock_nist_clock_sdram_controller_write2precharge_timer_count <= 3'd4;
		main_nist_clock_nist_clock_sdram_controller_refresh_timer_count <= 10'd975;
		main_nist_clock_nist_clock_adr_offset_r <= 4'd0;
		main_nist_clock_spiflash_bus_ack <= 1'd0;
		main_nist_clock_spiflash_bitbang_storage_full <= 4'd0;
		main_nist_clock_spiflash_bitbang_re <= 1'd0;
		main_nist_clock_spiflash_bitbang_en_storage_full <= 1'd0;
		main_nist_clock_spiflash_bitbang_en_re <= 1'd0;
		main_nist_clock_spiflash_cs_n1 <= 1'd1;
		main_nist_clock_spiflash_clk <= 1'd0;
		main_nist_clock_spiflash_dq_oe <= 1'd0;
		main_nist_clock_spiflash_sr <= 32'd0;
		main_nist_clock_spiflash_i1 <= 1'd0;
		main_nist_clock_spiflash_dqi <= 4'd0;
		main_nist_clock_spiflash_counter <= 7'd0;
		main_ethphy_mode0 <= 1'd0;
		main_ethphy_sys_counter <= 24'd0;
		main_ethphy_storage_full <= 1'd0;
		main_ethphy_re <= 1'd0;
		main_preamble_errors_status <= 32'd0;
		main_crc_errors_status <= 32'd0;
		main_tx_cdc_graycounter0_q <= 7'd0;
		main_tx_cdc_graycounter0_q_binary <= 7'd0;
		main_rx_cdc_graycounter1_q <= 7'd0;
		main_rx_cdc_graycounter1_q_binary <= 7'd0;
		main_writer_errors_status <= 32'd0;
		main_writer_storage_full <= 1'd0;
		main_writer_re <= 1'd0;
		main_writer_counter <= 32'd0;
		main_writer_slot <= 2'd0;
		main_writer_fifo_level <= 3'd0;
		main_writer_fifo_produce <= 2'd0;
		main_writer_fifo_consume <= 2'd0;
		main_reader_slot_storage_full <= 2'd0;
		main_reader_slot_re <= 1'd0;
		main_reader_length_storage_full <= 11'd0;
		main_reader_length_re <= 1'd0;
		main_reader_done_pending <= 1'd0;
		main_reader_eventmanager_storage_full <= 1'd0;
		main_reader_eventmanager_re <= 1'd0;
		main_reader_fifo_level <= 3'd0;
		main_reader_fifo_produce <= 2'd0;
		main_reader_fifo_consume <= 2'd0;
		main_reader_counter <= 11'd0;
		main_reader_last_d <= 1'd0;
		main_sram0_bus_ack0 <= 1'd0;
		main_sram1_bus_ack0 <= 1'd0;
		main_sram2_bus_ack0 <= 1'd0;
		main_sram3_bus_ack0 <= 1'd0;
		main_sram0_bus_ack1 <= 1'd0;
		main_sram1_bus_ack1 <= 1'd0;
		main_sram2_bus_ack1 <= 1'd0;
		main_sram3_bus_ack1 <= 1'd0;
		main_slave_sel_r <= 8'd0;
		main_kernel_cpu_storage_full <= 1'd1;
		main_kernel_cpu_re <= 1'd0;
		main_mailbox_i1_dat_r <= 32'd0;
		main_mailbox_i1_ack <= 1'd0;
		main_mailbox_i2_dat_r <= 32'd0;
		main_mailbox_i2_ack <= 1'd0;
		main_mailbox0 <= 32'd0;
		main_mailbox1 <= 32'd0;
		main_mailbox2 <= 32'd0;
		main_add_identifier_storage_full <= 8'd0;
		main_add_identifier_re <= 1'd0;
		main_load_storage_full <= 64'd0;
		main_load_re <= 1'd0;
		main_reload_storage_full <= 64'd0;
		main_reload_re <= 1'd0;
		main_en_storage_full <= 1'd0;
		main_en_re <= 1'd0;
		main_value_status <= 64'd0;
		main_zero_pending <= 1'd0;
		main_zero_old_trigger <= 1'd0;
		main_eventmanager_storage_full <= 1'd0;
		main_eventmanager_re <= 1'd0;
		main_value <= 64'd0;
		main_leds_storage_full <= 2'd0;
		main_leds_re <= 1'd0;
		main_i2c_out_storage_full <= 2'd0;
		main_i2c_out_re <= 1'd0;
		main_i2c_oe_storage_full <= 2'd0;
		main_i2c_oe_re <= 1'd0;
		main_rtio_crg_clock_sel_storage_full <= 1'd0;
		main_rtio_crg_clock_sel_re <= 1'd0;
		main_rtio_crg_pll_reset_storage_full <= 1'd1;
		main_rtio_crg_pll_reset_re <= 1'd0;
		main_rtio_core_collision_channel_status <= 16'd0;
		main_rtio_core_busy_channel_status <= 16'd0;
		main_rtio_core_sequence_error_channel_status <= 16'd0;
		main_rtio_core_cmd_reset <= 1'd1;
		main_rtio_core_cmd_reset_phy <= 1'd1;
		main_rtio_core_outputs_lanedistributor_minimum_coarse_timestamp <= 61'd0;
		main_rtio_core_o_collision <= 1'd0;
		main_rtio_core_o_busy <= 1'd0;
		main_rtio_core_o_sequence_error <= 1'd0;
		main_rtio_target_storage_full <= 32'd0;
		main_rtio_target_re <= 1'd0;
		main_rtio_o_data_storage_full <= 512'd0;
		main_rtio_o_data_re <= 1'd0;
		main_rtio_i_timeout_storage_full <= 64'd0;
		main_rtio_i_timeout_re <= 1'd0;
		main_rtio_counter_status <= 64'd0;
		main_rtio_now_hi_backing <= 32'd0;
		main_dma_dma_storage_full <= 36'd0;
		main_dma_dma_re <= 1'd0;
		main_dma_time_offset_storage_full <= 64'd0;
		main_dma_time_offset_re <= 1'd0;
		main_csrbank0_bus_dat_r <= 32'd0;
		main_csrbank0_bus_ack <= 1'd0;
		main_csrbank1_bus_dat_r <= 32'd0;
		main_csrbank1_bus_ack <= 1'd0;
		main_cri_con_storage_full <= 2'd0;
		main_cri_con_re <= 1'd0;
		main_cri_con_selected <= 1'd0;
		main_csrbank2_bus_dat_r <= 32'd0;
		main_csrbank2_bus_ack <= 1'd0;
		main_mon_chan_sel_storage_full <= 5'd0;
		main_mon_chan_sel_re <= 1'd0;
		main_mon_probe_sel_storage_full <= 4'd0;
		main_mon_probe_sel_re <= 1'd0;
		main_mon_status <= 32'd0;
		main_mon_bussynchronizer28_ping_o1 <= 1'd0;
		main_mon_bussynchronizer29_ping_o1 <= 1'd0;
		main_mon_bussynchronizer30_ping_o1 <= 1'd0;
		main_mon_bussynchronizer31_ping_o1 <= 1'd0;
		main_mon_bussynchronizer32_ping_o1 <= 1'd0;
		main_mon_bussynchronizer33_ping_o1 <= 1'd0;
		main_mon_bussynchronizer34_ping_o1 <= 1'd0;
		main_mon_bussynchronizer35_ping_o1 <= 1'd0;
		main_mon_bussynchronizer36_ping_o1 <= 1'd0;
		main_mon_bussynchronizer37_ping_o1 <= 1'd0;
		main_mon_bussynchronizer38_ping_o1 <= 1'd0;
		main_inj_chan_sel_storage_full <= 5'd0;
		main_inj_chan_sel_re <= 1'd0;
		main_inj_override_sel_storage_full <= 2'd0;
		main_inj_override_sel_re <= 1'd0;
		main_inj_o_sys0 <= 1'd0;
		main_inj_o_sys1 <= 1'd0;
		main_inj_o_sys2 <= 1'd0;
		main_inj_o_sys3 <= 1'd0;
		main_inj_o_sys4 <= 1'd0;
		main_inj_o_sys5 <= 1'd0;
		main_inj_o_sys6 <= 1'd0;
		main_inj_o_sys7 <= 1'd0;
		main_inj_o_sys8 <= 1'd0;
		main_inj_o_sys9 <= 1'd0;
		main_inj_o_sys10 <= 1'd0;
		main_inj_o_sys11 <= 1'd0;
		main_inj_o_sys12 <= 1'd0;
		main_inj_o_sys13 <= 1'd0;
		main_inj_o_sys14 <= 1'd0;
		main_inj_o_sys15 <= 1'd0;
		main_inj_o_sys16 <= 1'd0;
		main_inj_o_sys17 <= 1'd0;
		main_inj_o_sys18 <= 1'd0;
		main_inj_o_sys19 <= 1'd0;
		main_inj_o_sys20 <= 1'd0;
		main_inj_o_sys21 <= 1'd0;
		main_inj_o_sys22 <= 1'd0;
		main_inj_o_sys23 <= 1'd0;
		main_inj_o_sys24 <= 1'd0;
		main_inj_o_sys25 <= 1'd0;
		main_inj_o_sys26 <= 1'd0;
		main_inj_o_sys27 <= 1'd0;
		main_inj_o_sys28 <= 1'd0;
		main_inj_o_sys29 <= 1'd0;
		main_inj_o_sys30 <= 1'd0;
		main_inj_o_sys31 <= 1'd0;
		main_inj_o_sys32 <= 1'd0;
		main_inj_o_sys33 <= 1'd0;
		main_inj_o_sys34 <= 1'd0;
		main_inj_o_sys35 <= 1'd0;
		main_inj_o_sys36 <= 1'd0;
		main_inj_o_sys37 <= 1'd0;
		main_inj_o_sys38 <= 1'd0;
		main_inj_o_sys39 <= 1'd0;
		main_inj_o_sys40 <= 1'd0;
		main_inj_o_sys41 <= 1'd0;
		main_inj_o_sys42 <= 1'd0;
		main_inj_o_sys43 <= 1'd0;
		main_inj_o_sys44 <= 1'd0;
		main_inj_o_sys45 <= 1'd0;
		main_inj_o_sys46 <= 1'd0;
		main_inj_o_sys47 <= 1'd0;
		main_inj_o_sys48 <= 1'd0;
		main_interface1_bus_adr <= 30'd0;
		main_rtio_analyzer_enable_storage_full <= 1'd0;
		main_rtio_analyzer_enable_re <= 1'd0;
		main_rtio_analyzer_busy_status <= 1'd0;
		main_rtio_analyzer_message_encoder_source_stb <= 1'd0;
		main_rtio_analyzer_message_encoder_source_eop <= 1'd0;
		main_rtio_analyzer_message_encoder_source_payload_data <= 256'd0;
		main_rtio_analyzer_message_encoder_status <= 1'd0;
		main_rtio_analyzer_message_encoder_read_wait_event_r <= 1'd0;
		main_rtio_analyzer_message_encoder_just_written <= 1'd0;
		main_rtio_analyzer_message_encoder_enable_r <= 1'd0;
		main_rtio_analyzer_message_encoder_stopping <= 1'd0;
		main_rtio_analyzer_fifo_readable <= 1'd0;
		main_rtio_analyzer_fifo_level0 <= 8'd0;
		main_rtio_analyzer_fifo_produce <= 7'd0;
		main_rtio_analyzer_fifo_consume <= 7'd0;
		main_rtio_analyzer_converter_source_eop <= 1'd0;
		main_rtio_analyzer_converter_source_payload_data <= 512'd0;
		main_rtio_analyzer_converter_source_payload_valid_token_count <= 2'd0;
		main_rtio_analyzer_converter_demux <= 1'd0;
		main_rtio_analyzer_converter_strobe_all <= 1'd0;
		main_rtio_analyzer_dma_base_address_storage_full <= 36'd0;
		main_rtio_analyzer_dma_base_address_re <= 1'd0;
		main_rtio_analyzer_dma_last_address_storage_full <= 36'd0;
		main_rtio_analyzer_dma_last_address_re <= 1'd0;
		main_rtio_analyzer_dma_message_count <= 59'd0;
		main_rtio_analyzer_enable_r <= 1'd0;
		builder_minicon_state <= 5'd0;
		builder_fullmemorywe_state <= 3'd0;
		builder_liteethphygmiimii_state <= 2'd0;
		builder_liteethmacsramwriter_state <= 2'd0;
		builder_liteethmacsramreader_state <= 2'd0;
		builder_grant <= 1'd0;
		builder_slave_sel_r <= 5'd0;
		builder_sdram_cpulevel_arbiter_grant <= 1'd0;
		builder_sdram_native_arbiter_grant <= 2'd0;
		builder_nist_clock_grant <= 1'd0;
		builder_nist_clock_slave_sel_r <= 6'd0;
		builder_nist_clock_interface0_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface1_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface2_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface3_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface4_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface5_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface6_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface7_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface8_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface9_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface10_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface11_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface12_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface13_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface14_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface15_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface16_bank_bus_dat_r <= 8'd0;
		builder_nist_clock_interface17_bank_bus_dat_r <= 8'd0;
	end
	builder_xilinxmultiregimpl0_regs0 <= serial_rx;
	builder_xilinxmultiregimpl0_regs1 <= builder_xilinxmultiregimpl0_regs0;
	builder_xilinxmultiregimpl1_regs0 <= main_ethphy_toggle_i;
	builder_xilinxmultiregimpl1_regs1 <= builder_xilinxmultiregimpl1_regs0;
	builder_xilinxmultiregimpl2_regs0 <= main_ps_preamble_error_toggle_i;
	builder_xilinxmultiregimpl2_regs1 <= builder_xilinxmultiregimpl2_regs0;
	builder_xilinxmultiregimpl3_regs0 <= main_ps_crc_error_toggle_i;
	builder_xilinxmultiregimpl3_regs1 <= builder_xilinxmultiregimpl3_regs0;
	builder_xilinxmultiregimpl5_regs0 <= main_tx_cdc_graycounter1_q;
	builder_xilinxmultiregimpl5_regs1 <= builder_xilinxmultiregimpl5_regs0;
	builder_xilinxmultiregimpl6_regs0 <= main_rx_cdc_graycounter0_q;
	builder_xilinxmultiregimpl6_regs1 <= builder_xilinxmultiregimpl6_regs0;
	builder_xilinxmultiregimpl8_regs0 <= main_i2c_tstriple0_i;
	builder_xilinxmultiregimpl8_regs1 <= builder_xilinxmultiregimpl8_regs0;
	builder_xilinxmultiregimpl9_regs0 <= main_i2c_tstriple1_i;
	builder_xilinxmultiregimpl9_regs1 <= builder_xilinxmultiregimpl9_regs0;
	builder_xilinxmultiregimpl10_regs0 <= main_rtio_crg_pll_locked;
	builder_xilinxmultiregimpl10_regs1 <= builder_xilinxmultiregimpl10_regs0;
	builder_xilinxmultiregimpl11_regs0 <= main_value_gray_rtio;
	builder_xilinxmultiregimpl11_regs1 <= builder_xilinxmultiregimpl11_regs0;
	builder_xilinxmultiregimpl82_regs0 <= main_mon_bussynchronizer0_i;
	builder_xilinxmultiregimpl82_regs1 <= builder_xilinxmultiregimpl82_regs0;
	builder_xilinxmultiregimpl83_regs0 <= main_mon_bussynchronizer1_i;
	builder_xilinxmultiregimpl83_regs1 <= builder_xilinxmultiregimpl83_regs0;
	builder_xilinxmultiregimpl84_regs0 <= main_mon_bussynchronizer2_i;
	builder_xilinxmultiregimpl84_regs1 <= builder_xilinxmultiregimpl84_regs0;
	builder_xilinxmultiregimpl85_regs0 <= main_mon_bussynchronizer3_i;
	builder_xilinxmultiregimpl85_regs1 <= builder_xilinxmultiregimpl85_regs0;
	builder_xilinxmultiregimpl86_regs0 <= main_mon_bussynchronizer4_i;
	builder_xilinxmultiregimpl86_regs1 <= builder_xilinxmultiregimpl86_regs0;
	builder_xilinxmultiregimpl87_regs0 <= main_mon_bussynchronizer5_i;
	builder_xilinxmultiregimpl87_regs1 <= builder_xilinxmultiregimpl87_regs0;
	builder_xilinxmultiregimpl88_regs0 <= main_mon_bussynchronizer6_i;
	builder_xilinxmultiregimpl88_regs1 <= builder_xilinxmultiregimpl88_regs0;
	builder_xilinxmultiregimpl89_regs0 <= main_mon_bussynchronizer7_i;
	builder_xilinxmultiregimpl89_regs1 <= builder_xilinxmultiregimpl89_regs0;
	builder_xilinxmultiregimpl90_regs0 <= main_mon_bussynchronizer8_i;
	builder_xilinxmultiregimpl90_regs1 <= builder_xilinxmultiregimpl90_regs0;
	builder_xilinxmultiregimpl91_regs0 <= main_mon_bussynchronizer9_i;
	builder_xilinxmultiregimpl91_regs1 <= builder_xilinxmultiregimpl91_regs0;
	builder_xilinxmultiregimpl92_regs0 <= main_mon_bussynchronizer10_i;
	builder_xilinxmultiregimpl92_regs1 <= builder_xilinxmultiregimpl92_regs0;
	builder_xilinxmultiregimpl93_regs0 <= main_mon_bussynchronizer11_i;
	builder_xilinxmultiregimpl93_regs1 <= builder_xilinxmultiregimpl93_regs0;
	builder_xilinxmultiregimpl94_regs0 <= main_mon_bussynchronizer12_i;
	builder_xilinxmultiregimpl94_regs1 <= builder_xilinxmultiregimpl94_regs0;
	builder_xilinxmultiregimpl95_regs0 <= main_mon_bussynchronizer13_i;
	builder_xilinxmultiregimpl95_regs1 <= builder_xilinxmultiregimpl95_regs0;
	builder_xilinxmultiregimpl96_regs0 <= main_mon_bussynchronizer14_i;
	builder_xilinxmultiregimpl96_regs1 <= builder_xilinxmultiregimpl96_regs0;
	builder_xilinxmultiregimpl97_regs0 <= main_mon_bussynchronizer15_i;
	builder_xilinxmultiregimpl97_regs1 <= builder_xilinxmultiregimpl97_regs0;
	builder_xilinxmultiregimpl98_regs0 <= main_mon_bussynchronizer16_i;
	builder_xilinxmultiregimpl98_regs1 <= builder_xilinxmultiregimpl98_regs0;
	builder_xilinxmultiregimpl99_regs0 <= main_mon_bussynchronizer17_i;
	builder_xilinxmultiregimpl99_regs1 <= builder_xilinxmultiregimpl99_regs0;
	builder_xilinxmultiregimpl100_regs0 <= main_mon_bussynchronizer18_i;
	builder_xilinxmultiregimpl100_regs1 <= builder_xilinxmultiregimpl100_regs0;
	builder_xilinxmultiregimpl101_regs0 <= main_mon_bussynchronizer19_i;
	builder_xilinxmultiregimpl101_regs1 <= builder_xilinxmultiregimpl101_regs0;
	builder_xilinxmultiregimpl102_regs0 <= main_mon_bussynchronizer20_i;
	builder_xilinxmultiregimpl102_regs1 <= builder_xilinxmultiregimpl102_regs0;
	builder_xilinxmultiregimpl103_regs0 <= main_mon_bussynchronizer21_i;
	builder_xilinxmultiregimpl103_regs1 <= builder_xilinxmultiregimpl103_regs0;
	builder_xilinxmultiregimpl104_regs0 <= main_mon_bussynchronizer22_i;
	builder_xilinxmultiregimpl104_regs1 <= builder_xilinxmultiregimpl104_regs0;
	builder_xilinxmultiregimpl105_regs0 <= main_mon_bussynchronizer23_i;
	builder_xilinxmultiregimpl105_regs1 <= builder_xilinxmultiregimpl105_regs0;
	builder_xilinxmultiregimpl106_regs0 <= main_mon_bussynchronizer24_i;
	builder_xilinxmultiregimpl106_regs1 <= builder_xilinxmultiregimpl106_regs0;
	builder_xilinxmultiregimpl107_regs0 <= main_mon_bussynchronizer25_i;
	builder_xilinxmultiregimpl107_regs1 <= builder_xilinxmultiregimpl107_regs0;
	builder_xilinxmultiregimpl108_regs0 <= main_mon_bussynchronizer26_i;
	builder_xilinxmultiregimpl108_regs1 <= builder_xilinxmultiregimpl108_regs0;
	builder_xilinxmultiregimpl109_regs0 <= main_mon_bussynchronizer27_i;
	builder_xilinxmultiregimpl109_regs1 <= builder_xilinxmultiregimpl109_regs0;
	builder_xilinxmultiregimpl110_regs0 <= main_mon_bussynchronizer28_ping_toggle_i;
	builder_xilinxmultiregimpl110_regs1 <= builder_xilinxmultiregimpl110_regs0;
	builder_xilinxmultiregimpl112_regs0 <= main_mon_bussynchronizer28_ibuffer;
	builder_xilinxmultiregimpl112_regs1 <= builder_xilinxmultiregimpl112_regs0;
	builder_xilinxmultiregimpl113_regs0 <= main_mon_bussynchronizer29_ping_toggle_i;
	builder_xilinxmultiregimpl113_regs1 <= builder_xilinxmultiregimpl113_regs0;
	builder_xilinxmultiregimpl115_regs0 <= main_mon_bussynchronizer29_ibuffer;
	builder_xilinxmultiregimpl115_regs1 <= builder_xilinxmultiregimpl115_regs0;
	builder_xilinxmultiregimpl116_regs0 <= main_mon_bussynchronizer30_ping_toggle_i;
	builder_xilinxmultiregimpl116_regs1 <= builder_xilinxmultiregimpl116_regs0;
	builder_xilinxmultiregimpl118_regs0 <= main_mon_bussynchronizer30_ibuffer;
	builder_xilinxmultiregimpl118_regs1 <= builder_xilinxmultiregimpl118_regs0;
	builder_xilinxmultiregimpl119_regs0 <= main_mon_bussynchronizer31_ping_toggle_i;
	builder_xilinxmultiregimpl119_regs1 <= builder_xilinxmultiregimpl119_regs0;
	builder_xilinxmultiregimpl121_regs0 <= main_mon_bussynchronizer31_ibuffer;
	builder_xilinxmultiregimpl121_regs1 <= builder_xilinxmultiregimpl121_regs0;
	builder_xilinxmultiregimpl122_regs0 <= main_mon_bussynchronizer32_ping_toggle_i;
	builder_xilinxmultiregimpl122_regs1 <= builder_xilinxmultiregimpl122_regs0;
	builder_xilinxmultiregimpl124_regs0 <= main_mon_bussynchronizer32_ibuffer;
	builder_xilinxmultiregimpl124_regs1 <= builder_xilinxmultiregimpl124_regs0;
	builder_xilinxmultiregimpl125_regs0 <= main_mon_bussynchronizer33_ping_toggle_i;
	builder_xilinxmultiregimpl125_regs1 <= builder_xilinxmultiregimpl125_regs0;
	builder_xilinxmultiregimpl127_regs0 <= main_mon_bussynchronizer33_ibuffer;
	builder_xilinxmultiregimpl127_regs1 <= builder_xilinxmultiregimpl127_regs0;
	builder_xilinxmultiregimpl128_regs0 <= main_mon_bussynchronizer34_ping_toggle_i;
	builder_xilinxmultiregimpl128_regs1 <= builder_xilinxmultiregimpl128_regs0;
	builder_xilinxmultiregimpl130_regs0 <= main_mon_bussynchronizer34_ibuffer;
	builder_xilinxmultiregimpl130_regs1 <= builder_xilinxmultiregimpl130_regs0;
	builder_xilinxmultiregimpl131_regs0 <= main_mon_bussynchronizer35_ping_toggle_i;
	builder_xilinxmultiregimpl131_regs1 <= builder_xilinxmultiregimpl131_regs0;
	builder_xilinxmultiregimpl133_regs0 <= main_mon_bussynchronizer35_ibuffer;
	builder_xilinxmultiregimpl133_regs1 <= builder_xilinxmultiregimpl133_regs0;
	builder_xilinxmultiregimpl134_regs0 <= main_mon_bussynchronizer36_ping_toggle_i;
	builder_xilinxmultiregimpl134_regs1 <= builder_xilinxmultiregimpl134_regs0;
	builder_xilinxmultiregimpl136_regs0 <= main_mon_bussynchronizer36_ibuffer;
	builder_xilinxmultiregimpl136_regs1 <= builder_xilinxmultiregimpl136_regs0;
	builder_xilinxmultiregimpl137_regs0 <= main_mon_bussynchronizer37_ping_toggle_i;
	builder_xilinxmultiregimpl137_regs1 <= builder_xilinxmultiregimpl137_regs0;
	builder_xilinxmultiregimpl139_regs0 <= main_mon_bussynchronizer37_ibuffer;
	builder_xilinxmultiregimpl139_regs1 <= builder_xilinxmultiregimpl139_regs0;
	builder_xilinxmultiregimpl140_regs0 <= main_mon_bussynchronizer38_ping_toggle_i;
	builder_xilinxmultiregimpl140_regs1 <= builder_xilinxmultiregimpl140_regs0;
	builder_xilinxmultiregimpl142_regs0 <= main_mon_bussynchronizer38_ibuffer;
	builder_xilinxmultiregimpl142_regs1 <= builder_xilinxmultiregimpl142_regs0;
end

always @(posedge sys_kernel_clk) begin
	main_dma_dma_enable_r <= main_dma_flow_enable;
	if ((main_dma_flow_enable & (~main_dma_dma_enable_r))) begin
		main_dma_dma_sink_payload_address <= main_dma_dma_storage;
		main_dma_dma_sink_eop <= 1'd0;
		main_dma_dma_sink_stb <= 1'd1;
	end
	if ((main_dma_dma_sink_stb & main_dma_dma_sink_ack)) begin
		if (main_dma_dma_sink_eop) begin
			main_dma_dma_sink_stb <= 1'd0;
		end else begin
			main_dma_dma_sink_payload_address <= (main_dma_dma_sink_payload_address + 1'd1);
			if ((~main_dma_flow_enable)) begin
				main_dma_dma_sink_eop <= 1'd1;
			end
		end
	end
	if (main_dma_dma_source_ack) begin
		main_dma_dma_data_reg_loaded <= 1'd0;
	end
	if (main_interface0_bus_ack) begin
		main_dma_dma_data_reg_loaded <= 1'd1;
		main_dma_dma_source_payload_data <= main_interface0_bus_dat_r;
		main_dma_dma_source_eop <= main_dma_dma_sink_eop;
	end
	main_dma_rawslicer_level <= main_dma_rawslicer_next_level;
	if (main_dma_rawslicer_load_buf) begin
		case (main_dma_rawslicer_level)
			1'd0: begin
				main_dma_rawslicer_buf[511:0] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			1'd1: begin
				main_dma_rawslicer_buf[519:8] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			2'd2: begin
				main_dma_rawslicer_buf[527:16] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			2'd3: begin
				main_dma_rawslicer_buf[535:24] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			3'd4: begin
				main_dma_rawslicer_buf[543:32] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			3'd5: begin
				main_dma_rawslicer_buf[551:40] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			3'd6: begin
				main_dma_rawslicer_buf[559:48] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			3'd7: begin
				main_dma_rawslicer_buf[567:56] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd8: begin
				main_dma_rawslicer_buf[575:64] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd9: begin
				main_dma_rawslicer_buf[583:72] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd10: begin
				main_dma_rawslicer_buf[591:80] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd11: begin
				main_dma_rawslicer_buf[599:88] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd12: begin
				main_dma_rawslicer_buf[607:96] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd13: begin
				main_dma_rawslicer_buf[615:104] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd14: begin
				main_dma_rawslicer_buf[623:112] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			4'd15: begin
				main_dma_rawslicer_buf[631:120] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd16: begin
				main_dma_rawslicer_buf[639:128] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd17: begin
				main_dma_rawslicer_buf[647:136] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd18: begin
				main_dma_rawslicer_buf[655:144] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd19: begin
				main_dma_rawslicer_buf[663:152] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd20: begin
				main_dma_rawslicer_buf[671:160] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd21: begin
				main_dma_rawslicer_buf[679:168] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd22: begin
				main_dma_rawslicer_buf[687:176] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd23: begin
				main_dma_rawslicer_buf[695:184] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd24: begin
				main_dma_rawslicer_buf[703:192] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd25: begin
				main_dma_rawslicer_buf[711:200] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd26: begin
				main_dma_rawslicer_buf[719:208] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd27: begin
				main_dma_rawslicer_buf[727:216] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd28: begin
				main_dma_rawslicer_buf[735:224] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd29: begin
				main_dma_rawslicer_buf[743:232] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd30: begin
				main_dma_rawslicer_buf[751:240] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			5'd31: begin
				main_dma_rawslicer_buf[759:248] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd32: begin
				main_dma_rawslicer_buf[767:256] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd33: begin
				main_dma_rawslicer_buf[775:264] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd34: begin
				main_dma_rawslicer_buf[783:272] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd35: begin
				main_dma_rawslicer_buf[791:280] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd36: begin
				main_dma_rawslicer_buf[799:288] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd37: begin
				main_dma_rawslicer_buf[807:296] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd38: begin
				main_dma_rawslicer_buf[815:304] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd39: begin
				main_dma_rawslicer_buf[823:312] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd40: begin
				main_dma_rawslicer_buf[831:320] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd41: begin
				main_dma_rawslicer_buf[839:328] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd42: begin
				main_dma_rawslicer_buf[847:336] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd43: begin
				main_dma_rawslicer_buf[855:344] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd44: begin
				main_dma_rawslicer_buf[863:352] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd45: begin
				main_dma_rawslicer_buf[871:360] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd46: begin
				main_dma_rawslicer_buf[879:368] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd47: begin
				main_dma_rawslicer_buf[887:376] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd48: begin
				main_dma_rawslicer_buf[895:384] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd49: begin
				main_dma_rawslicer_buf[903:392] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd50: begin
				main_dma_rawslicer_buf[911:400] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd51: begin
				main_dma_rawslicer_buf[919:408] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd52: begin
				main_dma_rawslicer_buf[927:416] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd53: begin
				main_dma_rawslicer_buf[935:424] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd54: begin
				main_dma_rawslicer_buf[943:432] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd55: begin
				main_dma_rawslicer_buf[951:440] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd56: begin
				main_dma_rawslicer_buf[959:448] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd57: begin
				main_dma_rawslicer_buf[967:456] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd58: begin
				main_dma_rawslicer_buf[975:464] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd59: begin
				main_dma_rawslicer_buf[983:472] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd60: begin
				main_dma_rawslicer_buf[991:480] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd61: begin
				main_dma_rawslicer_buf[999:488] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd62: begin
				main_dma_rawslicer_buf[1007:496] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			6'd63: begin
				main_dma_rawslicer_buf[1015:504] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd64: begin
				main_dma_rawslicer_buf[1023:512] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd65: begin
				main_dma_rawslicer_buf[1031:520] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd66: begin
				main_dma_rawslicer_buf[1039:528] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd67: begin
				main_dma_rawslicer_buf[1047:536] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd68: begin
				main_dma_rawslicer_buf[1055:544] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd69: begin
				main_dma_rawslicer_buf[1063:552] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd70: begin
				main_dma_rawslicer_buf[1071:560] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd71: begin
				main_dma_rawslicer_buf[1079:568] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd72: begin
				main_dma_rawslicer_buf[1087:576] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd73: begin
				main_dma_rawslicer_buf[1095:584] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd74: begin
				main_dma_rawslicer_buf[1103:592] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd75: begin
				main_dma_rawslicer_buf[1111:600] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
			7'd76: begin
				main_dma_rawslicer_buf[1119:608] <= {main_dma_rawslicer_sink_payload_data[7:0], main_dma_rawslicer_sink_payload_data[15:8], main_dma_rawslicer_sink_payload_data[23:16], main_dma_rawslicer_sink_payload_data[31:24], main_dma_rawslicer_sink_payload_data[39:32], main_dma_rawslicer_sink_payload_data[47:40], main_dma_rawslicer_sink_payload_data[55:48], main_dma_rawslicer_sink_payload_data[63:56], main_dma_rawslicer_sink_payload_data[71:64], main_dma_rawslicer_sink_payload_data[79:72], main_dma_rawslicer_sink_payload_data[87:80], main_dma_rawslicer_sink_payload_data[95:88], main_dma_rawslicer_sink_payload_data[103:96], main_dma_rawslicer_sink_payload_data[111:104], main_dma_rawslicer_sink_payload_data[119:112], main_dma_rawslicer_sink_payload_data[127:120], main_dma_rawslicer_sink_payload_data[135:128], main_dma_rawslicer_sink_payload_data[143:136], main_dma_rawslicer_sink_payload_data[151:144], main_dma_rawslicer_sink_payload_data[159:152], main_dma_rawslicer_sink_payload_data[167:160], main_dma_rawslicer_sink_payload_data[175:168], main_dma_rawslicer_sink_payload_data[183:176], main_dma_rawslicer_sink_payload_data[191:184], main_dma_rawslicer_sink_payload_data[199:192], main_dma_rawslicer_sink_payload_data[207:200], main_dma_rawslicer_sink_payload_data[215:208], main_dma_rawslicer_sink_payload_data[223:216], main_dma_rawslicer_sink_payload_data[231:224], main_dma_rawslicer_sink_payload_data[239:232], main_dma_rawslicer_sink_payload_data[247:240], main_dma_rawslicer_sink_payload_data[255:248], main_dma_rawslicer_sink_payload_data[263:256], main_dma_rawslicer_sink_payload_data[271:264], main_dma_rawslicer_sink_payload_data[279:272], main_dma_rawslicer_sink_payload_data[287:280], main_dma_rawslicer_sink_payload_data[295:288], main_dma_rawslicer_sink_payload_data[303:296], main_dma_rawslicer_sink_payload_data[311:304], main_dma_rawslicer_sink_payload_data[319:312], main_dma_rawslicer_sink_payload_data[327:320], main_dma_rawslicer_sink_payload_data[335:328], main_dma_rawslicer_sink_payload_data[343:336], main_dma_rawslicer_sink_payload_data[351:344], main_dma_rawslicer_sink_payload_data[359:352], main_dma_rawslicer_sink_payload_data[367:360], main_dma_rawslicer_sink_payload_data[375:368], main_dma_rawslicer_sink_payload_data[383:376], main_dma_rawslicer_sink_payload_data[391:384], main_dma_rawslicer_sink_payload_data[399:392], main_dma_rawslicer_sink_payload_data[407:400], main_dma_rawslicer_sink_payload_data[415:408], main_dma_rawslicer_sink_payload_data[423:416], main_dma_rawslicer_sink_payload_data[431:424], main_dma_rawslicer_sink_payload_data[439:432], main_dma_rawslicer_sink_payload_data[447:440], main_dma_rawslicer_sink_payload_data[455:448], main_dma_rawslicer_sink_payload_data[463:456], main_dma_rawslicer_sink_payload_data[471:464], main_dma_rawslicer_sink_payload_data[479:472], main_dma_rawslicer_sink_payload_data[487:480], main_dma_rawslicer_sink_payload_data[495:488], main_dma_rawslicer_sink_payload_data[503:496], main_dma_rawslicer_sink_payload_data[511:504]};
			end
		endcase
	end
	if (main_dma_rawslicer_shift_buf) begin
		case (main_dma_rawslicer_source_consume)
			1'd0: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:0];
			end
			1'd1: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:8];
			end
			2'd2: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:16];
			end
			2'd3: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:24];
			end
			3'd4: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:32];
			end
			3'd5: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:40];
			end
			3'd6: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:48];
			end
			3'd7: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:56];
			end
			4'd8: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:64];
			end
			4'd9: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:72];
			end
			4'd10: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:80];
			end
			4'd11: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:88];
			end
			4'd12: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:96];
			end
			4'd13: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:104];
			end
			4'd14: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:112];
			end
			4'd15: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:120];
			end
			5'd16: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:128];
			end
			5'd17: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:136];
			end
			5'd18: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:144];
			end
			5'd19: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:152];
			end
			5'd20: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:160];
			end
			5'd21: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:168];
			end
			5'd22: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:176];
			end
			5'd23: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:184];
			end
			5'd24: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:192];
			end
			5'd25: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:200];
			end
			5'd26: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:208];
			end
			5'd27: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:216];
			end
			5'd28: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:224];
			end
			5'd29: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:232];
			end
			5'd30: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:240];
			end
			5'd31: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:248];
			end
			6'd32: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:256];
			end
			6'd33: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:264];
			end
			6'd34: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:272];
			end
			6'd35: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:280];
			end
			6'd36: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:288];
			end
			6'd37: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:296];
			end
			6'd38: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:304];
			end
			6'd39: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:312];
			end
			6'd40: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:320];
			end
			6'd41: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:328];
			end
			6'd42: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:336];
			end
			6'd43: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:344];
			end
			6'd44: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:352];
			end
			6'd45: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:360];
			end
			6'd46: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:368];
			end
			6'd47: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:376];
			end
			6'd48: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:384];
			end
			6'd49: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:392];
			end
			6'd50: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:400];
			end
			6'd51: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:408];
			end
			6'd52: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:416];
			end
			6'd53: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:424];
			end
			6'd54: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:432];
			end
			6'd55: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:440];
			end
			6'd56: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:448];
			end
			6'd57: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:456];
			end
			6'd58: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:464];
			end
			6'd59: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:472];
			end
			6'd60: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:480];
			end
			6'd61: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:488];
			end
			6'd62: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:496];
			end
			6'd63: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:504];
			end
			7'd64: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:512];
			end
			7'd65: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:520];
			end
			7'd66: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:528];
			end
			7'd67: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:536];
			end
			7'd68: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:544];
			end
			7'd69: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:552];
			end
			7'd70: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:560];
			end
			7'd71: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:568];
			end
			7'd72: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:576];
			end
			7'd73: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:584];
			end
			7'd74: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:592];
			end
			7'd75: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:600];
			end
			7'd76: begin
				main_dma_rawslicer_buf <= main_dma_rawslicer_buf[1119:608];
			end
		endcase
	end
	builder_resetinserter_state <= builder_resetinserter_next_state;
	if (main_dma_reset) begin
		main_dma_rawslicer_buf <= 1120'd0;
		main_dma_rawslicer_level <= 8'd0;
		builder_resetinserter_state <= 2'd0;
	end
	builder_recordconverter_state <= builder_recordconverter_next_state;
	if (main_dma_time_offset_source_ack) begin
		main_dma_time_offset_source_stb <= 1'd0;
	end
	if ((~main_dma_time_offset_source_stb)) begin
		main_dma_time_offset_source_payload_length <= main_dma_time_offset_sink_payload_length;
		main_dma_time_offset_source_payload_channel <= main_dma_time_offset_sink_payload_channel;
		main_dma_time_offset_source_payload_address <= main_dma_time_offset_sink_payload_address;
		main_dma_time_offset_source_payload_data <= main_dma_time_offset_sink_payload_data;
		main_dma_time_offset_source_payload_timestamp <= (main_dma_time_offset_sink_payload_timestamp + main_dma_time_offset_storage);
		main_dma_time_offset_source_eop <= main_dma_time_offset_sink_eop;
		main_dma_time_offset_source_stb <= main_dma_time_offset_sink_stb;
	end
	if (main_dma_cri_master_underflow_trigger) begin
		main_dma_cri_master_error_w <= 1'd1;
		main_dma_cri_master_error_channel_status <= main_dma_cri_master_sink_payload_channel;
		main_dma_cri_master_error_timestamp_status <= main_dma_cri_master_sink_payload_timestamp;
		main_dma_cri_master_error_address_status <= main_dma_cri_master_sink_payload_address;
	end
	if (main_dma_cri_master_link_error_trigger) begin
		main_dma_cri_master_error_w <= 2'd2;
		main_dma_cri_master_error_channel_status <= main_dma_cri_master_sink_payload_channel;
		main_dma_cri_master_error_timestamp_status <= main_dma_cri_master_sink_payload_timestamp;
		main_dma_cri_master_error_address_status <= main_dma_cri_master_sink_payload_address;
	end
	if (main_dma_cri_master_error_re) begin
		main_dma_cri_master_error_w <= 1'd0;
	end
	builder_crimaster_state <= builder_crimaster_next_state;
	builder_fsm_state <= builder_fsm_next_state;
	if (sys_kernel_rst) begin
		main_dma_dma_sink_stb <= 1'd0;
		main_dma_dma_sink_eop <= 1'd0;
		main_dma_dma_sink_payload_address <= 30'd0;
		main_dma_dma_source_eop <= 1'd0;
		main_dma_dma_source_payload_data <= 512'd0;
		main_dma_dma_data_reg_loaded <= 1'd0;
		main_dma_dma_enable_r <= 1'd0;
		main_dma_rawslicer_buf <= 1120'd0;
		main_dma_rawslicer_level <= 8'd0;
		main_dma_time_offset_source_stb <= 1'd0;
		main_dma_time_offset_source_eop <= 1'd0;
		main_dma_time_offset_source_payload_length <= 8'd0;
		main_dma_time_offset_source_payload_channel <= 24'd0;
		main_dma_time_offset_source_payload_timestamp <= 64'd0;
		main_dma_time_offset_source_payload_address <= 8'd0;
		main_dma_time_offset_source_payload_data <= 512'd0;
		main_dma_cri_master_error_w <= 2'd0;
		main_dma_cri_master_error_channel_status <= 24'd0;
		main_dma_cri_master_error_timestamp_status <= 64'd0;
		main_dma_cri_master_error_address_status <= 16'd0;
		builder_resetinserter_state <= 2'd0;
		builder_recordconverter_state <= 2'd0;
		builder_crimaster_state <= 3'd0;
		builder_fsm_state <= 3'd0;
	end
end

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(24'd11468800)
) mor1kx (
	.clk(sys_clk),
	.dwbm_ack_i(main_nist_clock_nist_clock_dbus_ack),
	.dwbm_dat_i(main_nist_clock_nist_clock_dbus_dat_r),
	.dwbm_err_i(main_nist_clock_nist_clock_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(main_nist_clock_nist_clock_interrupt),
	.iwbm_ack_i(main_nist_clock_nist_clock_ibus_ack),
	.iwbm_dat_i(main_nist_clock_nist_clock_ibus_dat_r),
	.iwbm_err_i(main_nist_clock_nist_clock_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_rst),
	.dwbm_adr_o(main_nist_clock_nist_clock_d_adr_o),
	.dwbm_bte_o(main_nist_clock_nist_clock_dbus_bte),
	.dwbm_cti_o(main_nist_clock_nist_clock_dbus_cti),
	.dwbm_cyc_o(main_nist_clock_nist_clock_dbus_cyc),
	.dwbm_dat_o(main_nist_clock_nist_clock_dbus_dat_w),
	.dwbm_sel_o(main_nist_clock_nist_clock_dbus_sel),
	.dwbm_stb_o(main_nist_clock_nist_clock_dbus_stb),
	.dwbm_we_o(main_nist_clock_nist_clock_dbus_we),
	.iwbm_adr_o(main_nist_clock_nist_clock_i_adr_o),
	.iwbm_bte_o(main_nist_clock_nist_clock_ibus_bte),
	.iwbm_cti_o(main_nist_clock_nist_clock_ibus_cti),
	.iwbm_cyc_o(main_nist_clock_nist_clock_ibus_cyc),
	.iwbm_dat_o(main_nist_clock_nist_clock_ibus_dat_w),
	.iwbm_sel_o(main_nist_clock_nist_clock_ibus_sel),
	.iwbm_stb_o(main_nist_clock_nist_clock_ibus_stb),
	.iwbm_we_o(main_nist_clock_nist_clock_ibus_we)
);

reg [31:0] mem[0:2047];
reg [10:0] memadr;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_sram_we[0])
		mem[main_nist_clock_nist_clock_sram_adr][7:0] <= main_nist_clock_nist_clock_sram_dat_w[7:0];
	if (main_nist_clock_nist_clock_sram_we[1])
		mem[main_nist_clock_nist_clock_sram_adr][15:8] <= main_nist_clock_nist_clock_sram_dat_w[15:8];
	if (main_nist_clock_nist_clock_sram_we[2])
		mem[main_nist_clock_nist_clock_sram_adr][23:16] <= main_nist_clock_nist_clock_sram_dat_w[23:16];
	if (main_nist_clock_nist_clock_sram_we[3])
		mem[main_nist_clock_nist_clock_sram_adr][31:24] <= main_nist_clock_nist_clock_sram_dat_w[31:24];
	memadr <= main_nist_clock_nist_clock_sram_adr;
end

assign main_nist_clock_nist_clock_sram_dat_r = mem[memadr];

reg [8:0] storage[0:15];
reg [8:0] memdat;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_uart_tx_fifo_wrport_we)
		storage[main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr] <= main_nist_clock_nist_clock_uart_tx_fifo_wrport_dat_w;
	memdat <= storage[main_nist_clock_nist_clock_uart_tx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_nist_clock_nist_clock_uart_tx_fifo_wrport_dat_r = memdat;
assign main_nist_clock_nist_clock_uart_tx_fifo_rdport_dat_r = storage[main_nist_clock_nist_clock_uart_tx_fifo_rdport_adr];

reg [8:0] storage_1[0:15];
reg [8:0] memdat_1;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_uart_rx_fifo_wrport_we)
		storage_1[main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr] <= main_nist_clock_nist_clock_uart_rx_fifo_wrport_dat_w;
	memdat_1 <= storage_1[main_nist_clock_nist_clock_uart_rx_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_nist_clock_nist_clock_uart_rx_fifo_wrport_dat_r = memdat_1;
assign main_nist_clock_nist_clock_uart_rx_fifo_rdport_dat_r = storage_1[main_nist_clock_nist_clock_uart_rx_fifo_rdport_adr];

IBUFDS IBUFDS(
	.I(clk200_p),
	.IB(clk200_n),
	.O(main_nist_clock_clk200_se)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(3'd5),
	.CLKIN1_PERIOD(5.0),
	.CLKOUT0_DIVIDE(4'd8),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(3'd5),
	.CLKOUT2_PHASE(0.0),
	.CLKOUT3_DIVIDE(2'd2),
	.CLKOUT3_PHASE(0.0),
	.CLKOUT4_DIVIDE(3'd4),
	.CLKOUT4_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE (
	.CLKFBIN(main_nist_clock_pll_fb),
	.CLKIN1(main_nist_clock_clk200_se),
	.CLKFBOUT(main_nist_clock_pll_fb),
	.CLKOUT0(main_nist_clock_pll_sys),
	.CLKOUT1(main_nist_clock_pll_sys4x),
	.CLKOUT2(main_nist_clock_pll_clk200),
	.LOCKED(main_nist_clock_pll_locked)
);

BUFG BUFG(
	.I(main_nist_clock_pll_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(main_nist_clock_pll_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_2(
	.I(main_nist_clock_pll_clk200),
	.O(clk200_clk)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(main_nist_clock_ic_reset)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(main_nist_clock_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[0]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[0]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[0]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[0]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[0]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[0]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[0]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[1]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[1]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[1]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[1]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[1]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[1]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[1]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[2]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[2]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[2]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[2]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[2]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[2]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[2]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[3]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[3]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[3]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[3]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[3]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[3]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[3]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[4]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[4]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[4]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[4]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[4]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[4]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[4]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[5]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[5]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[5]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[5]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[5]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[5]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[5]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[6]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[6]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[6]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[6]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[6]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[6]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[6]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[7]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[7]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[7]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[7]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[7]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[7]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[7]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[8]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[8]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[8]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[8]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[8]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[8]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[8]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[9]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[9]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[9]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[9]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[9]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[9]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[9]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[10]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[10]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[10]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[10]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[10]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[10]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[10]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[11]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[11]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[11]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[11]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[11]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[11]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[11]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[12]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[12]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[12]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[12]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[12]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[12]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[12]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[13]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[13]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[13]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[13]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[13]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[13]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[13]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[14]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[14]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[14]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[14]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[14]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[14]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[14]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_address[15]),
	.D2(main_nist_clock_ddrphy_dfi_p0_address[15]),
	.D3(main_nist_clock_ddrphy_dfi_p1_address[15]),
	.D4(main_nist_clock_ddrphy_dfi_p1_address[15]),
	.D5(main_nist_clock_ddrphy_dfi_p2_address[15]),
	.D6(main_nist_clock_ddrphy_dfi_p2_address[15]),
	.D7(main_nist_clock_ddrphy_dfi_p3_address[15]),
	.D8(main_nist_clock_ddrphy_dfi_p3_address[15]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[15])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_bank[0]),
	.D2(main_nist_clock_ddrphy_dfi_p0_bank[0]),
	.D3(main_nist_clock_ddrphy_dfi_p1_bank[0]),
	.D4(main_nist_clock_ddrphy_dfi_p1_bank[0]),
	.D5(main_nist_clock_ddrphy_dfi_p2_bank[0]),
	.D6(main_nist_clock_ddrphy_dfi_p2_bank[0]),
	.D7(main_nist_clock_ddrphy_dfi_p3_bank[0]),
	.D8(main_nist_clock_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_bank[1]),
	.D2(main_nist_clock_ddrphy_dfi_p0_bank[1]),
	.D3(main_nist_clock_ddrphy_dfi_p1_bank[1]),
	.D4(main_nist_clock_ddrphy_dfi_p1_bank[1]),
	.D5(main_nist_clock_ddrphy_dfi_p2_bank[1]),
	.D6(main_nist_clock_ddrphy_dfi_p2_bank[1]),
	.D7(main_nist_clock_ddrphy_dfi_p3_bank[1]),
	.D8(main_nist_clock_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_bank[2]),
	.D2(main_nist_clock_ddrphy_dfi_p0_bank[2]),
	.D3(main_nist_clock_ddrphy_dfi_p1_bank[2]),
	.D4(main_nist_clock_ddrphy_dfi_p1_bank[2]),
	.D5(main_nist_clock_ddrphy_dfi_p2_bank[2]),
	.D6(main_nist_clock_ddrphy_dfi_p2_bank[2]),
	.D7(main_nist_clock_ddrphy_dfi_p3_bank[2]),
	.D8(main_nist_clock_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_ras_n),
	.D2(main_nist_clock_ddrphy_dfi_p0_ras_n),
	.D3(main_nist_clock_ddrphy_dfi_p1_ras_n),
	.D4(main_nist_clock_ddrphy_dfi_p1_ras_n),
	.D5(main_nist_clock_ddrphy_dfi_p2_ras_n),
	.D6(main_nist_clock_ddrphy_dfi_p2_ras_n),
	.D7(main_nist_clock_ddrphy_dfi_p3_ras_n),
	.D8(main_nist_clock_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_cas_n),
	.D2(main_nist_clock_ddrphy_dfi_p0_cas_n),
	.D3(main_nist_clock_ddrphy_dfi_p1_cas_n),
	.D4(main_nist_clock_ddrphy_dfi_p1_cas_n),
	.D5(main_nist_clock_ddrphy_dfi_p2_cas_n),
	.D6(main_nist_clock_ddrphy_dfi_p2_cas_n),
	.D7(main_nist_clock_ddrphy_dfi_p3_cas_n),
	.D8(main_nist_clock_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_we_n),
	.D2(main_nist_clock_ddrphy_dfi_p0_we_n),
	.D3(main_nist_clock_ddrphy_dfi_p1_we_n),
	.D4(main_nist_clock_ddrphy_dfi_p1_we_n),
	.D5(main_nist_clock_ddrphy_dfi_p2_we_n),
	.D6(main_nist_clock_ddrphy_dfi_p2_we_n),
	.D7(main_nist_clock_ddrphy_dfi_p3_we_n),
	.D8(main_nist_clock_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_cs_n),
	.D2(main_nist_clock_ddrphy_dfi_p0_cs_n),
	.D3(main_nist_clock_ddrphy_dfi_p1_cs_n),
	.D4(main_nist_clock_ddrphy_dfi_p1_cs_n),
	.D5(main_nist_clock_ddrphy_dfi_p2_cs_n),
	.D6(main_nist_clock_ddrphy_dfi_p2_cs_n),
	.D7(main_nist_clock_ddrphy_dfi_p3_cs_n),
	.D8(main_nist_clock_ddrphy_dfi_p3_cs_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cs_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_cke),
	.D2(main_nist_clock_ddrphy_dfi_p0_cke),
	.D3(main_nist_clock_ddrphy_dfi_p1_cke),
	.D4(main_nist_clock_ddrphy_dfi_p1_cke),
	.D5(main_nist_clock_ddrphy_dfi_p2_cke),
	.D6(main_nist_clock_ddrphy_dfi_p2_cke),
	.D7(main_nist_clock_ddrphy_dfi_p3_cke),
	.D8(main_nist_clock_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_odt),
	.D2(main_nist_clock_ddrphy_dfi_p0_odt),
	.D3(main_nist_clock_ddrphy_dfi_p1_odt),
	.D4(main_nist_clock_ddrphy_dfi_p1_odt),
	.D5(main_nist_clock_ddrphy_dfi_p2_odt),
	.D6(main_nist_clock_ddrphy_dfi_p2_odt),
	.D7(main_nist_clock_ddrphy_dfi_p3_odt),
	.D8(main_nist_clock_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_reset_n),
	.D2(main_nist_clock_ddrphy_dfi_p0_reset_n),
	.D3(main_nist_clock_ddrphy_dfi_p1_reset_n),
	.D4(main_nist_clock_ddrphy_dfi_p1_reset_n),
	.D5(main_nist_clock_ddrphy_dfi_p2_reset_n),
	.D6(main_nist_clock_ddrphy_dfi_p2_reset_n),
	.D7(main_nist_clock_ddrphy_dfi_p3_reset_n),
	.D8(main_nist_clock_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[8]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[8]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[8]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay0)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[0]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay0),
	.TQ(main_nist_clock_ddrphy_dqs_t0)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_1 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed0),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay0)
);

OBUFTDS OBUFTDS(
	.I(main_nist_clock_ddrphy_dqs_delayed0),
	.T(main_nist_clock_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[9]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[9]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[9]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay1)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_2 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[1]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay1),
	.TQ(main_nist_clock_ddrphy_dqs_t1)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_3 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed1),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay1)
);

OBUFTDS OBUFTDS_1(
	.I(main_nist_clock_ddrphy_dqs_delayed1),
	.T(main_nist_clock_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[2]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[10]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[2]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[10]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[2]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[10]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[2]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay2)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_4 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[2]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay2),
	.TQ(main_nist_clock_ddrphy_dqs_t2)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_5 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed2),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay2)
);

OBUFTDS OBUFTDS_2(
	.I(main_nist_clock_ddrphy_dqs_delayed2),
	.T(main_nist_clock_ddrphy_dqs_t2),
	.O(ddram_dqs_p[2]),
	.OB(ddram_dqs_n[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[3]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[11]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[3]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[11]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[3]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[11]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[3]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay3)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_6 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[3]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay3),
	.TQ(main_nist_clock_ddrphy_dqs_t3)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_7 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed3),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay3)
);

OBUFTDS OBUFTDS_3(
	.I(main_nist_clock_ddrphy_dqs_delayed3),
	.T(main_nist_clock_ddrphy_dqs_t3),
	.O(ddram_dqs_p[3]),
	.OB(ddram_dqs_n[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[4]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[12]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[4]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[12]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[4]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[12]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[4]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay4)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_8 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[4]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay4),
	.TQ(main_nist_clock_ddrphy_dqs_t4)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_9 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed4),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay4)
);

OBUFTDS OBUFTDS_4(
	.I(main_nist_clock_ddrphy_dqs_delayed4),
	.T(main_nist_clock_ddrphy_dqs_t4),
	.O(ddram_dqs_p[4]),
	.OB(ddram_dqs_n[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[5]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[13]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[5]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[13]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[5]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[13]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[5]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay5)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_10 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[5]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay5),
	.TQ(main_nist_clock_ddrphy_dqs_t5)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_11 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed5),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay5)
);

OBUFTDS OBUFTDS_5(
	.I(main_nist_clock_ddrphy_dqs_delayed5),
	.T(main_nist_clock_ddrphy_dqs_t5),
	.O(ddram_dqs_p[5]),
	.OB(ddram_dqs_n[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[6]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[14]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[6]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[14]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[6]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[14]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[6]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay6)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_12 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[6]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay6),
	.TQ(main_nist_clock_ddrphy_dqs_t6)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_13 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed6),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay6)
);

OBUFTDS OBUFTDS_6(
	.I(main_nist_clock_ddrphy_dqs_delayed6),
	.T(main_nist_clock_ddrphy_dqs_t6),
	.O(ddram_dqs_p[6]),
	.OB(ddram_dqs_n[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[7]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata_mask[15]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[7]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata_mask[15]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[7]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata_mask[15]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[7]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata_mask[15]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_nist_clock_ddrphy_dm_o_nodelay7)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_14 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(ddram_dm[7]),
	.ODATAIN(main_nist_clock_ddrphy_dm_o_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dqs_serdes_pattern[0]),
	.D2(main_nist_clock_ddrphy_dqs_serdes_pattern[1]),
	.D3(main_nist_clock_ddrphy_dqs_serdes_pattern[2]),
	.D4(main_nist_clock_ddrphy_dqs_serdes_pattern[3]),
	.D5(main_nist_clock_ddrphy_dqs_serdes_pattern[4]),
	.D6(main_nist_clock_ddrphy_dqs_serdes_pattern[5]),
	.D7(main_nist_clock_ddrphy_dqs_serdes_pattern[6]),
	.D8(main_nist_clock_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_nist_clock_ddrphy_dqs_nodelay7),
	.TQ(main_nist_clock_ddrphy_dqs_t7)
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_15 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dqs_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dqs_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dqs_delayed7),
	.ODATAIN(main_nist_clock_ddrphy_dqs_nodelay7)
);

OBUFTDS OBUFTDS_7(
	.I(main_nist_clock_ddrphy_dqs_delayed7),
	.T(main_nist_clock_ddrphy_dqs_t7),
	.O(ddram_dqs_p[7]),
	.OB(ddram_dqs_n[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[0]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[64]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[0]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[64]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[0]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[64]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[0]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[64]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay0),
	.TQ(main_nist_clock_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[64]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[0]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[64]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[0]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[64]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[0]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[64]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[0])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_16 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed0),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay0)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(main_nist_clock_ddrphy_dq_o_delayed0),
	.T(main_nist_clock_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[1]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[65]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[1]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[65]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[1]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[65]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[1]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[65]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay1),
	.TQ(main_nist_clock_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[65]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[1]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[65]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[1]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[65]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[1]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[65]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[1])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_17 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed1),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay1)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(main_nist_clock_ddrphy_dq_o_delayed1),
	.T(main_nist_clock_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[2]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[66]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[2]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[66]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[2]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[66]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[2]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[66]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay2),
	.TQ(main_nist_clock_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[66]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[2]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[66]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[2]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[66]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[2]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[66]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[2])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_18 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed2),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay2)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(main_nist_clock_ddrphy_dq_o_delayed2),
	.T(main_nist_clock_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[3]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[67]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[3]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[67]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[3]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[67]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[3]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[67]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay3),
	.TQ(main_nist_clock_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[67]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[3]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[67]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[3]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[67]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[3]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[67]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[3])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_19 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed3),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay3)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(main_nist_clock_ddrphy_dq_o_delayed3),
	.T(main_nist_clock_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[4]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[68]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[4]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[68]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[4]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[68]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[4]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[68]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay4),
	.TQ(main_nist_clock_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[68]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[4]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[68]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[4]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[68]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[4]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[68]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[4])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_20 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed4),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay4)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(main_nist_clock_ddrphy_dq_o_delayed4),
	.T(main_nist_clock_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[5]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[69]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[5]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[69]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[5]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[69]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[5]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[69]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay5),
	.TQ(main_nist_clock_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[69]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[5]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[69]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[5]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[69]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[5]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[69]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[5])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_21 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed5),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay5)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(main_nist_clock_ddrphy_dq_o_delayed5),
	.T(main_nist_clock_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[6]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[70]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[6]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[70]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[6]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[70]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[6]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[70]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay6),
	.TQ(main_nist_clock_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[70]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[6]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[70]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[6]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[70]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[6]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[70]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[6])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_22 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed6),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay6)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(main_nist_clock_ddrphy_dq_o_delayed6),
	.T(main_nist_clock_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[7]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[71]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[7]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[71]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[7]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[71]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[7]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[71]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay7),
	.TQ(main_nist_clock_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[71]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[7]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[71]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[7]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[71]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[7]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[71]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[7])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_23 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed7),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay7)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[0] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(main_nist_clock_ddrphy_dq_o_delayed7),
	.T(main_nist_clock_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[8]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[72]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[8]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[72]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[8]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[72]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[8]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[72]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay8),
	.TQ(main_nist_clock_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[72]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[8]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[72]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[8]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[72]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[8]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[72]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[8])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_24 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed8),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay8)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(main_nist_clock_ddrphy_dq_o_delayed8),
	.T(main_nist_clock_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[9]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[73]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[9]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[73]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[9]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[73]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[9]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[73]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay9),
	.TQ(main_nist_clock_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[73]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[9]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[73]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[9]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[73]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[9]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[73]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[9])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_25 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed9),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay9)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(main_nist_clock_ddrphy_dq_o_delayed9),
	.T(main_nist_clock_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_53 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[10]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[74]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[10]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[74]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[10]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[74]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[10]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[74]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay10),
	.TQ(main_nist_clock_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[74]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[10]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[74]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[10]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[74]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[10]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[74]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[10])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_26 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed10),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay10)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(main_nist_clock_ddrphy_dq_o_delayed10),
	.T(main_nist_clock_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_54 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[11]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[75]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[11]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[75]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[11]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[75]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[11]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[75]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay11),
	.TQ(main_nist_clock_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[75]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[11]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[75]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[11]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[75]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[11]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[75]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[11])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_27 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed11),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay11)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(main_nist_clock_ddrphy_dq_o_delayed11),
	.T(main_nist_clock_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_55 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[12]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[76]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[12]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[76]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[12]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[76]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[12]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[76]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay12),
	.TQ(main_nist_clock_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[76]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[12]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[76]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[12]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[76]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[12]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[76]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[12])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_28 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed12),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay12)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(main_nist_clock_ddrphy_dq_o_delayed12),
	.T(main_nist_clock_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_56 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[13]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[77]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[13]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[77]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[13]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[77]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[13]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[77]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay13),
	.TQ(main_nist_clock_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[77]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[13]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[77]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[13]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[77]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[13]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[77]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[13])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_29 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed13),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay13)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(main_nist_clock_ddrphy_dq_o_delayed13),
	.T(main_nist_clock_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_57 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[14]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[78]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[14]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[78]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[14]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[78]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[14]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[78]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay14),
	.TQ(main_nist_clock_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[78]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[14]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[78]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[14]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[78]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[14]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[78]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[14])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_30 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed14),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay14)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(main_nist_clock_ddrphy_dq_o_delayed14),
	.T(main_nist_clock_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_58 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[15]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[79]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[15]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[79]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[15]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[79]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[15]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[79]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay15),
	.TQ(main_nist_clock_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[79]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[15]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[79]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[15]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[79]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[15]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[79]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[15])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_31 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed15),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay15)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[1] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(main_nist_clock_ddrphy_dq_o_delayed15),
	.T(main_nist_clock_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay15)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_59 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[16]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[80]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[16]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[80]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[16]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[80]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[16]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[80]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay16),
	.TQ(main_nist_clock_ddrphy_dq_t16)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_16 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed16),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[80]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[16]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[80]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[16]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[80]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[16]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[80]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[16])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_32 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed16),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay16)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_16 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay16),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed16)
);

IOBUF IOBUF_16(
	.I(main_nist_clock_ddrphy_dq_o_delayed16),
	.T(main_nist_clock_ddrphy_dq_t16),
	.IO(ddram_dq[16]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay16)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_60 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[17]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[81]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[17]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[81]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[17]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[81]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[17]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[81]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay17),
	.TQ(main_nist_clock_ddrphy_dq_t17)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_17 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed17),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[81]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[17]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[81]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[17]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[81]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[17]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[81]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[17])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_33 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed17),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay17)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_17 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay17),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed17)
);

IOBUF IOBUF_17(
	.I(main_nist_clock_ddrphy_dq_o_delayed17),
	.T(main_nist_clock_ddrphy_dq_t17),
	.IO(ddram_dq[17]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay17)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_61 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[18]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[82]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[18]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[82]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[18]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[82]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[18]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[82]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay18),
	.TQ(main_nist_clock_ddrphy_dq_t18)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_18 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed18),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[82]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[18]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[82]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[18]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[82]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[18]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[82]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[18])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_34 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed18),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay18)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_18 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay18),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed18)
);

IOBUF IOBUF_18(
	.I(main_nist_clock_ddrphy_dq_o_delayed18),
	.T(main_nist_clock_ddrphy_dq_t18),
	.IO(ddram_dq[18]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay18)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_62 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[19]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[83]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[19]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[83]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[19]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[83]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[19]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[83]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay19),
	.TQ(main_nist_clock_ddrphy_dq_t19)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_19 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed19),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[83]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[19]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[83]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[19]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[83]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[19]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[83]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[19])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_35 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed19),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay19)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_19 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay19),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed19)
);

IOBUF IOBUF_19(
	.I(main_nist_clock_ddrphy_dq_o_delayed19),
	.T(main_nist_clock_ddrphy_dq_t19),
	.IO(ddram_dq[19]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay19)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_63 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[20]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[84]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[20]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[84]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[20]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[84]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[20]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[84]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay20),
	.TQ(main_nist_clock_ddrphy_dq_t20)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_20 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed20),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[84]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[20]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[84]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[20]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[84]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[20]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[84]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[20])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_36 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed20),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay20)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_20 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay20),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed20)
);

IOBUF IOBUF_20(
	.I(main_nist_clock_ddrphy_dq_o_delayed20),
	.T(main_nist_clock_ddrphy_dq_t20),
	.IO(ddram_dq[20]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay20)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_64 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[21]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[85]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[21]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[85]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[21]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[85]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[21]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[85]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay21),
	.TQ(main_nist_clock_ddrphy_dq_t21)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_21 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed21),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[85]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[21]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[85]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[21]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[85]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[21]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[85]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[21])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_37 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed21),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay21)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_21 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay21),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed21)
);

IOBUF IOBUF_21(
	.I(main_nist_clock_ddrphy_dq_o_delayed21),
	.T(main_nist_clock_ddrphy_dq_t21),
	.IO(ddram_dq[21]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay21)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_65 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[22]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[86]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[22]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[86]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[22]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[86]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[22]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[86]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay22),
	.TQ(main_nist_clock_ddrphy_dq_t22)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_22 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed22),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[86]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[22]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[86]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[22]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[86]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[22]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[86]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[22])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_38 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed22),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay22)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_22 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay22),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed22)
);

IOBUF IOBUF_22(
	.I(main_nist_clock_ddrphy_dq_o_delayed22),
	.T(main_nist_clock_ddrphy_dq_t22),
	.IO(ddram_dq[22]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay22)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_66 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[23]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[87]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[23]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[87]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[23]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[87]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[23]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[87]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay23),
	.TQ(main_nist_clock_ddrphy_dq_t23)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_23 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed23),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[87]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[23]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[87]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[23]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[87]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[23]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[87]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[23])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_39 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed23),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay23)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_23 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay23),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[2] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed23)
);

IOBUF IOBUF_23(
	.I(main_nist_clock_ddrphy_dq_o_delayed23),
	.T(main_nist_clock_ddrphy_dq_t23),
	.IO(ddram_dq[23]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay23)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_67 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[24]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[88]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[24]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[88]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[24]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[88]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[24]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[88]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay24),
	.TQ(main_nist_clock_ddrphy_dq_t24)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_24 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed24),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[88]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[24]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[88]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[24]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[88]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[24]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[88]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[24])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_40 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed24),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay24)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_24 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay24),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed24)
);

IOBUF IOBUF_24(
	.I(main_nist_clock_ddrphy_dq_o_delayed24),
	.T(main_nist_clock_ddrphy_dq_t24),
	.IO(ddram_dq[24]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay24)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_68 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[25]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[89]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[25]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[89]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[25]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[89]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[25]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[89]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay25),
	.TQ(main_nist_clock_ddrphy_dq_t25)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_25 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed25),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[89]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[25]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[89]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[25]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[89]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[25]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[89]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[25])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_41 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed25),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay25)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_25 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay25),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed25)
);

IOBUF IOBUF_25(
	.I(main_nist_clock_ddrphy_dq_o_delayed25),
	.T(main_nist_clock_ddrphy_dq_t25),
	.IO(ddram_dq[25]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay25)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_69 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[26]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[90]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[26]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[90]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[26]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[90]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[26]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[90]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay26),
	.TQ(main_nist_clock_ddrphy_dq_t26)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_26 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed26),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[90]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[26]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[90]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[26]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[90]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[26]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[90]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[26])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_42 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed26),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay26)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_26 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay26),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed26)
);

IOBUF IOBUF_26(
	.I(main_nist_clock_ddrphy_dq_o_delayed26),
	.T(main_nist_clock_ddrphy_dq_t26),
	.IO(ddram_dq[26]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay26)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_70 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[27]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[91]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[27]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[91]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[27]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[91]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[27]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[91]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay27),
	.TQ(main_nist_clock_ddrphy_dq_t27)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_27 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed27),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[91]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[27]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[91]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[27]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[91]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[27]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[91]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[27])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_43 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed27),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay27)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_27 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay27),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed27)
);

IOBUF IOBUF_27(
	.I(main_nist_clock_ddrphy_dq_o_delayed27),
	.T(main_nist_clock_ddrphy_dq_t27),
	.IO(ddram_dq[27]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay27)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_71 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[28]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[92]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[28]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[92]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[28]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[92]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[28]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[92]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay28),
	.TQ(main_nist_clock_ddrphy_dq_t28)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_28 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed28),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[92]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[28]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[92]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[28]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[92]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[28]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[92]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[28])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_44 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed28),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay28)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_28 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay28),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed28)
);

IOBUF IOBUF_28(
	.I(main_nist_clock_ddrphy_dq_o_delayed28),
	.T(main_nist_clock_ddrphy_dq_t28),
	.IO(ddram_dq[28]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay28)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_72 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[29]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[93]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[29]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[93]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[29]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[93]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[29]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[93]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay29),
	.TQ(main_nist_clock_ddrphy_dq_t29)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_29 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed29),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[93]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[29]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[93]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[29]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[93]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[29]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[93]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[29])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_45 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed29),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay29)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_29 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay29),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed29)
);

IOBUF IOBUF_29(
	.I(main_nist_clock_ddrphy_dq_o_delayed29),
	.T(main_nist_clock_ddrphy_dq_t29),
	.IO(ddram_dq[29]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay29)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_73 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[30]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[94]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[30]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[94]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[30]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[94]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[30]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[94]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay30),
	.TQ(main_nist_clock_ddrphy_dq_t30)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_30 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed30),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[94]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[30]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[94]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[30]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[94]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[30]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[94]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[30])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_46 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed30),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay30)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_30 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay30),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed30)
);

IOBUF IOBUF_30(
	.I(main_nist_clock_ddrphy_dq_o_delayed30),
	.T(main_nist_clock_ddrphy_dq_t30),
	.IO(ddram_dq[30]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay30)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_74 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[31]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[95]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[31]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[95]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[31]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[95]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[31]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[95]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay31),
	.TQ(main_nist_clock_ddrphy_dq_t31)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_31 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed31),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[95]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[31]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[95]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[31]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[95]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[31]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[95]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[31])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_47 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed31),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay31)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_31 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay31),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[3] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed31)
);

IOBUF IOBUF_31(
	.I(main_nist_clock_ddrphy_dq_o_delayed31),
	.T(main_nist_clock_ddrphy_dq_t31),
	.IO(ddram_dq[31]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay31)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_75 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[32]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[96]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[32]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[96]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[32]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[96]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[32]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[96]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay32),
	.TQ(main_nist_clock_ddrphy_dq_t32)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_32 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed32),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[96]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[32]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[96]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[32]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[96]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[32]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[96]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[32])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_48 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed32),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay32)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_32 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay32),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed32)
);

IOBUF IOBUF_32(
	.I(main_nist_clock_ddrphy_dq_o_delayed32),
	.T(main_nist_clock_ddrphy_dq_t32),
	.IO(ddram_dq[32]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay32)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_76 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[33]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[97]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[33]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[97]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[33]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[97]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[33]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[97]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay33),
	.TQ(main_nist_clock_ddrphy_dq_t33)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_33 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed33),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[97]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[33]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[97]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[33]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[97]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[33]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[97]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[33])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_49 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed33),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay33)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_33 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay33),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed33)
);

IOBUF IOBUF_33(
	.I(main_nist_clock_ddrphy_dq_o_delayed33),
	.T(main_nist_clock_ddrphy_dq_t33),
	.IO(ddram_dq[33]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay33)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_77 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[34]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[98]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[34]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[98]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[34]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[98]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[34]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[98]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay34),
	.TQ(main_nist_clock_ddrphy_dq_t34)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_34 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed34),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[98]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[34]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[98]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[34]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[98]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[34]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[98]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[34])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_50 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed34),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay34)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_34 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay34),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed34)
);

IOBUF IOBUF_34(
	.I(main_nist_clock_ddrphy_dq_o_delayed34),
	.T(main_nist_clock_ddrphy_dq_t34),
	.IO(ddram_dq[34]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay34)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_78 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[35]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[99]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[35]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[99]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[35]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[99]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[35]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[99]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay35),
	.TQ(main_nist_clock_ddrphy_dq_t35)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_35 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed35),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[99]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[35]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[99]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[35]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[99]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[35]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[99]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[35])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_51 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed35),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay35)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_35 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay35),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed35)
);

IOBUF IOBUF_35(
	.I(main_nist_clock_ddrphy_dq_o_delayed35),
	.T(main_nist_clock_ddrphy_dq_t35),
	.IO(ddram_dq[35]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay35)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_79 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[36]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[100]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[36]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[100]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[36]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[100]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[36]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[100]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay36),
	.TQ(main_nist_clock_ddrphy_dq_t36)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_36 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed36),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[100]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[36]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[100]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[36]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[100]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[36]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[100]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[36])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_52 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed36),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay36)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_36 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay36),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed36)
);

IOBUF IOBUF_36(
	.I(main_nist_clock_ddrphy_dq_o_delayed36),
	.T(main_nist_clock_ddrphy_dq_t36),
	.IO(ddram_dq[36]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay36)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_80 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[37]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[101]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[37]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[101]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[37]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[101]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[37]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[101]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay37),
	.TQ(main_nist_clock_ddrphy_dq_t37)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_37 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed37),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[101]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[37]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[101]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[37]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[101]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[37]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[101]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[37])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_53 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed37),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay37)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_37 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay37),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed37)
);

IOBUF IOBUF_37(
	.I(main_nist_clock_ddrphy_dq_o_delayed37),
	.T(main_nist_clock_ddrphy_dq_t37),
	.IO(ddram_dq[37]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay37)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_81 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[38]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[102]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[38]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[102]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[38]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[102]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[38]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[102]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay38),
	.TQ(main_nist_clock_ddrphy_dq_t38)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_38 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed38),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[102]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[38]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[102]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[38]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[102]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[38]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[102]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[38])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_54 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed38),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay38)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_38 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay38),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed38)
);

IOBUF IOBUF_38(
	.I(main_nist_clock_ddrphy_dq_o_delayed38),
	.T(main_nist_clock_ddrphy_dq_t38),
	.IO(ddram_dq[38]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay38)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_82 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[39]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[103]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[39]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[103]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[39]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[103]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[39]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[103]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay39),
	.TQ(main_nist_clock_ddrphy_dq_t39)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_39 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed39),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[103]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[39]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[103]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[39]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[103]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[39]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[103]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[39])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_55 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed39),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay39)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_39 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay39),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[4] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed39)
);

IOBUF IOBUF_39(
	.I(main_nist_clock_ddrphy_dq_o_delayed39),
	.T(main_nist_clock_ddrphy_dq_t39),
	.IO(ddram_dq[39]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay39)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_83 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[40]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[104]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[40]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[104]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[40]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[104]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[40]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[104]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay40),
	.TQ(main_nist_clock_ddrphy_dq_t40)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_40 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed40),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[104]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[40]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[104]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[40]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[104]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[40]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[104]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[40])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_56 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed40),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay40)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_40 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay40),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed40)
);

IOBUF IOBUF_40(
	.I(main_nist_clock_ddrphy_dq_o_delayed40),
	.T(main_nist_clock_ddrphy_dq_t40),
	.IO(ddram_dq[40]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay40)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_84 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[41]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[105]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[41]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[105]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[41]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[105]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[41]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[105]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay41),
	.TQ(main_nist_clock_ddrphy_dq_t41)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_41 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed41),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[105]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[41]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[105]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[41]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[105]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[41]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[105]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[41])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_57 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed41),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay41)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_41 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay41),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed41)
);

IOBUF IOBUF_41(
	.I(main_nist_clock_ddrphy_dq_o_delayed41),
	.T(main_nist_clock_ddrphy_dq_t41),
	.IO(ddram_dq[41]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay41)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_85 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[42]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[106]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[42]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[106]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[42]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[106]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[42]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[106]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay42),
	.TQ(main_nist_clock_ddrphy_dq_t42)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_42 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed42),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[106]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[42]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[106]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[42]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[106]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[42]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[106]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[42])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_58 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed42),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay42)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_42 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay42),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed42)
);

IOBUF IOBUF_42(
	.I(main_nist_clock_ddrphy_dq_o_delayed42),
	.T(main_nist_clock_ddrphy_dq_t42),
	.IO(ddram_dq[42]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay42)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_86 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[43]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[107]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[43]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[107]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[43]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[107]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[43]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[107]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay43),
	.TQ(main_nist_clock_ddrphy_dq_t43)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_43 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed43),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[107]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[43]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[107]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[43]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[107]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[43]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[107]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[43])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_59 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed43),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay43)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_43 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay43),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed43)
);

IOBUF IOBUF_43(
	.I(main_nist_clock_ddrphy_dq_o_delayed43),
	.T(main_nist_clock_ddrphy_dq_t43),
	.IO(ddram_dq[43]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay43)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_87 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[44]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[108]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[44]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[108]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[44]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[108]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[44]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[108]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay44),
	.TQ(main_nist_clock_ddrphy_dq_t44)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_44 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed44),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[108]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[44]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[108]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[44]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[108]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[44]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[108]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[44])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_60 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed44),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay44)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_44 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay44),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed44)
);

IOBUF IOBUF_44(
	.I(main_nist_clock_ddrphy_dq_o_delayed44),
	.T(main_nist_clock_ddrphy_dq_t44),
	.IO(ddram_dq[44]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay44)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_88 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[45]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[109]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[45]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[109]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[45]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[109]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[45]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[109]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay45),
	.TQ(main_nist_clock_ddrphy_dq_t45)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_45 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed45),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[109]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[45]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[109]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[45]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[109]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[45]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[109]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[45])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_61 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed45),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay45)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_45 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay45),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed45)
);

IOBUF IOBUF_45(
	.I(main_nist_clock_ddrphy_dq_o_delayed45),
	.T(main_nist_clock_ddrphy_dq_t45),
	.IO(ddram_dq[45]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay45)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_89 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[46]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[110]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[46]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[110]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[46]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[110]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[46]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[110]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay46),
	.TQ(main_nist_clock_ddrphy_dq_t46)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_46 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed46),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[110]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[46]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[110]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[46]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[110]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[46]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[110]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[46])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_62 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed46),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay46)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_46 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay46),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed46)
);

IOBUF IOBUF_46(
	.I(main_nist_clock_ddrphy_dq_o_delayed46),
	.T(main_nist_clock_ddrphy_dq_t46),
	.IO(ddram_dq[46]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay46)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_90 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[47]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[111]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[47]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[111]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[47]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[111]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[47]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[111]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay47),
	.TQ(main_nist_clock_ddrphy_dq_t47)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_47 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed47),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[111]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[47]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[111]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[47]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[111]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[47]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[111]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[47])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_63 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed47),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay47)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_47 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay47),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[5] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed47)
);

IOBUF IOBUF_47(
	.I(main_nist_clock_ddrphy_dq_o_delayed47),
	.T(main_nist_clock_ddrphy_dq_t47),
	.IO(ddram_dq[47]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay47)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_91 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[48]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[112]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[48]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[112]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[48]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[112]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[48]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[112]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay48),
	.TQ(main_nist_clock_ddrphy_dq_t48)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_48 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed48),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[112]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[48]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[112]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[48]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[112]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[48]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[112]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[48])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_64 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed48),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay48)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_48 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay48),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed48)
);

IOBUF IOBUF_48(
	.I(main_nist_clock_ddrphy_dq_o_delayed48),
	.T(main_nist_clock_ddrphy_dq_t48),
	.IO(ddram_dq[48]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay48)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_92 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[49]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[113]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[49]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[113]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[49]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[113]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[49]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[113]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay49),
	.TQ(main_nist_clock_ddrphy_dq_t49)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_49 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed49),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[113]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[49]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[113]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[49]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[113]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[49]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[113]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[49])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_65 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed49),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay49)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_49 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay49),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed49)
);

IOBUF IOBUF_49(
	.I(main_nist_clock_ddrphy_dq_o_delayed49),
	.T(main_nist_clock_ddrphy_dq_t49),
	.IO(ddram_dq[49]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay49)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_93 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[50]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[114]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[50]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[114]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[50]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[114]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[50]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[114]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay50),
	.TQ(main_nist_clock_ddrphy_dq_t50)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_50 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed50),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[114]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[50]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[114]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[50]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[114]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[50]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[114]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[50])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_66 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed50),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay50)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_50 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay50),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed50)
);

IOBUF IOBUF_50(
	.I(main_nist_clock_ddrphy_dq_o_delayed50),
	.T(main_nist_clock_ddrphy_dq_t50),
	.IO(ddram_dq[50]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay50)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_94 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[51]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[115]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[51]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[115]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[51]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[115]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[51]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[115]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay51),
	.TQ(main_nist_clock_ddrphy_dq_t51)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_51 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed51),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[115]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[51]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[115]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[51]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[115]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[51]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[115]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[51])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_67 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed51),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay51)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_51 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay51),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed51)
);

IOBUF IOBUF_51(
	.I(main_nist_clock_ddrphy_dq_o_delayed51),
	.T(main_nist_clock_ddrphy_dq_t51),
	.IO(ddram_dq[51]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay51)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_95 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[52]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[116]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[52]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[116]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[52]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[116]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[52]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[116]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay52),
	.TQ(main_nist_clock_ddrphy_dq_t52)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_52 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed52),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[116]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[52]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[116]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[52]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[116]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[52]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[116]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[52])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_68 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed52),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay52)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_52 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay52),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed52)
);

IOBUF IOBUF_52(
	.I(main_nist_clock_ddrphy_dq_o_delayed52),
	.T(main_nist_clock_ddrphy_dq_t52),
	.IO(ddram_dq[52]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay52)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_96 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[53]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[117]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[53]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[117]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[53]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[117]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[53]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[117]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay53),
	.TQ(main_nist_clock_ddrphy_dq_t53)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_53 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed53),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[117]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[53]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[117]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[53]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[117]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[53]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[117]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[53])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_69 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed53),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay53)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_53 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay53),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed53)
);

IOBUF IOBUF_53(
	.I(main_nist_clock_ddrphy_dq_o_delayed53),
	.T(main_nist_clock_ddrphy_dq_t53),
	.IO(ddram_dq[53]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay53)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_97 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[54]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[118]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[54]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[118]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[54]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[118]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[54]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[118]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay54),
	.TQ(main_nist_clock_ddrphy_dq_t54)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_54 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed54),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[118]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[54]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[118]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[54]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[118]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[54]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[118]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[54])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_70 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed54),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay54)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_54 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay54),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed54)
);

IOBUF IOBUF_54(
	.I(main_nist_clock_ddrphy_dq_o_delayed54),
	.T(main_nist_clock_ddrphy_dq_t54),
	.IO(ddram_dq[54]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay54)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_98 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[55]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[119]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[55]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[119]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[55]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[119]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[55]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[119]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay55),
	.TQ(main_nist_clock_ddrphy_dq_t55)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_55 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed55),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[119]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[55]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[119]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[55]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[119]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[55]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[119]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[55])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_71 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed55),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay55)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_55 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay55),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[6] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed55)
);

IOBUF IOBUF_55(
	.I(main_nist_clock_ddrphy_dq_o_delayed55),
	.T(main_nist_clock_ddrphy_dq_t55),
	.IO(ddram_dq[55]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay55)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_99 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[56]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[120]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[56]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[120]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[56]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[120]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[56]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[120]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay56),
	.TQ(main_nist_clock_ddrphy_dq_t56)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_56 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed56),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[120]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[56]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[120]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[56]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[120]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[56]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[120]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[56])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_72 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed56),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay56)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_56 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay56),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed56)
);

IOBUF IOBUF_56(
	.I(main_nist_clock_ddrphy_dq_o_delayed56),
	.T(main_nist_clock_ddrphy_dq_t56),
	.IO(ddram_dq[56]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay56)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_100 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[57]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[121]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[57]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[121]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[57]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[121]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[57]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[121]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay57),
	.TQ(main_nist_clock_ddrphy_dq_t57)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_57 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed57),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[121]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[57]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[121]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[57]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[121]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[57]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[121]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[57])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_73 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed57),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay57)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_57 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay57),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed57)
);

IOBUF IOBUF_57(
	.I(main_nist_clock_ddrphy_dq_o_delayed57),
	.T(main_nist_clock_ddrphy_dq_t57),
	.IO(ddram_dq[57]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay57)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_101 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[58]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[122]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[58]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[122]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[58]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[122]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[58]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[122]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay58),
	.TQ(main_nist_clock_ddrphy_dq_t58)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_58 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed58),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[122]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[58]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[122]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[58]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[122]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[58]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[122]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[58])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_74 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed58),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay58)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_58 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay58),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed58)
);

IOBUF IOBUF_58(
	.I(main_nist_clock_ddrphy_dq_o_delayed58),
	.T(main_nist_clock_ddrphy_dq_t58),
	.IO(ddram_dq[58]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay58)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_102 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[59]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[123]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[59]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[123]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[59]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[123]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[59]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[123]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay59),
	.TQ(main_nist_clock_ddrphy_dq_t59)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_59 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed59),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[123]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[59]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[123]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[59]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[123]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[59]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[123]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[59])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_75 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed59),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay59)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_59 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay59),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed59)
);

IOBUF IOBUF_59(
	.I(main_nist_clock_ddrphy_dq_o_delayed59),
	.T(main_nist_clock_ddrphy_dq_t59),
	.IO(ddram_dq[59]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay59)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_103 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[60]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[124]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[60]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[124]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[60]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[124]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[60]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[124]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay60),
	.TQ(main_nist_clock_ddrphy_dq_t60)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_60 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed60),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[124]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[60]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[124]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[60]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[124]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[60]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[124]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[60])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_76 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed60),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay60)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_60 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay60),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed60)
);

IOBUF IOBUF_60(
	.I(main_nist_clock_ddrphy_dq_o_delayed60),
	.T(main_nist_clock_ddrphy_dq_t60),
	.IO(ddram_dq[60]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay60)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_104 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[61]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[125]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[61]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[125]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[61]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[125]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[61]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[125]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay61),
	.TQ(main_nist_clock_ddrphy_dq_t61)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_61 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed61),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[125]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[61]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[125]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[61]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[125]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[61]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[125]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[61])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_77 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed61),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay61)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_61 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay61),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed61)
);

IOBUF IOBUF_61(
	.I(main_nist_clock_ddrphy_dq_o_delayed61),
	.T(main_nist_clock_ddrphy_dq_t61),
	.IO(ddram_dq[61]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay61)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_105 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[62]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[126]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[62]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[126]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[62]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[126]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[62]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[126]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay62),
	.TQ(main_nist_clock_ddrphy_dq_t62)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_62 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed62),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[126]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[62]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[126]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[62]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[126]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[62]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[126]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[62])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_78 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed62),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay62)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_62 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay62),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed62)
);

IOBUF IOBUF_62(
	.I(main_nist_clock_ddrphy_dq_o_delayed62),
	.T(main_nist_clock_ddrphy_dq_t62),
	.IO(ddram_dq[62]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay62)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_106 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_nist_clock_ddrphy_dfi_p0_wrdata[63]),
	.D2(main_nist_clock_ddrphy_dfi_p0_wrdata[127]),
	.D3(main_nist_clock_ddrphy_dfi_p1_wrdata[63]),
	.D4(main_nist_clock_ddrphy_dfi_p1_wrdata[127]),
	.D5(main_nist_clock_ddrphy_dfi_p2_wrdata[63]),
	.D6(main_nist_clock_ddrphy_dfi_p2_wrdata[127]),
	.D7(main_nist_clock_ddrphy_dfi_p3_wrdata[63]),
	.D8(main_nist_clock_ddrphy_dfi_p3_wrdata[127]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_nist_clock_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_nist_clock_ddrphy_dq_o_nodelay63),
	.TQ(main_nist_clock_ddrphy_dq_t63)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_63 (
	.BITSLIP((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(main_nist_clock_ddrphy_dq_i_delayed63),
	.RST((sys_rst | (main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re))),
	.Q1(main_nist_clock_ddrphy_dfi_p3_rddata[127]),
	.Q2(main_nist_clock_ddrphy_dfi_p3_rddata[63]),
	.Q3(main_nist_clock_ddrphy_dfi_p2_rddata[127]),
	.Q4(main_nist_clock_ddrphy_dfi_p2_rddata[63]),
	.Q5(main_nist_clock_ddrphy_dfi_p1_rddata[127]),
	.Q6(main_nist_clock_ddrphy_dfi_p1_rddata[63]),
	.Q7(main_nist_clock_ddrphy_dfi_p0_rddata[127]),
	.Q8(main_nist_clock_ddrphy_dfi_p0_rddata[63])
);

ODELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("ODATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.ODELAY_TYPE("VARIABLE"),
	.ODELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) ODELAYE2_79 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_inc_re)),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_wdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_o_delayed63),
	.ODATAIN(main_nist_clock_ddrphy_dq_o_nodelay63)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_63 (
	.C(sys_clk),
	.CE((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_nist_clock_ddrphy_dq_i_nodelay63),
	.INC(1'd1),
	.LD((main_nist_clock_ddrphy_dly_sel_storage[7] & main_nist_clock_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_nist_clock_ddrphy_dq_i_delayed63)
);

IOBUF IOBUF_63(
	.I(main_nist_clock_ddrphy_dq_o_delayed63),
	.T(main_nist_clock_ddrphy_dq_t63),
	.IO(ddram_dq[63]),
	.O(main_nist_clock_ddrphy_dq_i_nodelay63)
);

reg [23:0] tag_mem[0:2047];
reg [10:0] memadr_1;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_tag_port_we)
		tag_mem[main_nist_clock_nist_clock_tag_port_adr] <= main_nist_clock_nist_clock_tag_port_dat_w;
	memadr_1 <= main_nist_clock_nist_clock_tag_port_adr;
end

assign main_nist_clock_nist_clock_tag_port_dat_r = tag_mem[memadr_1];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(main_nist_clock_clk),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

assign spiflash_dq = main_nist_clock_spiflash_oe ? main_nist_clock_spiflash_o : 4'bz;
assign main_nist_clock_spiflash_i0 = spiflash_dq;

BUFGMUX BUFGMUX(
	.I0(eth_rx_clk),
	.I1(eth_clocks_tx),
	.S((main_ethphy_mode0 == 1'd1)),
	.O(eth_tx_clk)
);

reg [10:0] storage_2[0:4];
reg [10:0] memdat_2;
always @(posedge eth_rx_clk) begin
	if (main_crc32_checker_syncfifo_wrport_we)
		storage_2[main_crc32_checker_syncfifo_wrport_adr] <= main_crc32_checker_syncfifo_wrport_dat_w;
	memdat_2 <= storage_2[main_crc32_checker_syncfifo_wrport_adr];
end

always @(posedge eth_rx_clk) begin
end

assign main_crc32_checker_syncfifo_wrport_dat_r = memdat_2;
assign main_crc32_checker_syncfifo_rdport_dat_r = storage_2[main_crc32_checker_syncfifo_rdport_adr];

reg [40:0] storage_3[0:63];
reg [5:0] memadr_2;
reg [5:0] memadr_3;
always @(posedge sys_clk) begin
	if (main_tx_cdc_wrport_we)
		storage_3[main_tx_cdc_wrport_adr] <= main_tx_cdc_wrport_dat_w;
	memadr_2 <= main_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memadr_3 <= main_tx_cdc_rdport_adr;
end

assign main_tx_cdc_wrport_dat_r = storage_3[memadr_2];
assign main_tx_cdc_rdport_dat_r = storage_3[memadr_3];

reg [40:0] storage_4[0:63];
reg [5:0] memadr_4;
reg [5:0] memadr_5;
always @(posedge eth_rx_clk) begin
	if (main_rx_cdc_wrport_we)
		storage_4[main_rx_cdc_wrport_adr] <= main_rx_cdc_wrport_dat_w;
	memadr_4 <= main_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin
	memadr_5 <= main_rx_cdc_rdport_adr;
end

assign main_rx_cdc_wrport_dat_r = storage_4[memadr_4];
assign main_rx_cdc_rdport_dat_r = storage_4[memadr_5];

reg [34:0] storage_5[0:3];
reg [34:0] memdat_3;
always @(posedge sys_clk) begin
	if (main_writer_fifo_wrport_we)
		storage_5[main_writer_fifo_wrport_adr] <= main_writer_fifo_wrport_dat_w;
	memdat_3 <= storage_5[main_writer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_writer_fifo_wrport_dat_r = memdat_3;
assign main_writer_fifo_rdport_dat_r = storage_5[main_writer_fifo_rdport_adr];

reg [31:0] mem_1[0:381];
reg [8:0] memadr_6;
reg [8:0] memadr_7;
always @(posedge sys_clk) begin
	if (main_writer_memory0_we)
		mem_1[main_writer_memory0_adr] <= main_writer_memory0_dat_w;
	memadr_6 <= main_writer_memory0_adr;
end

always @(posedge sys_clk) begin
	memadr_7 <= main_sram0_adr0;
end

assign main_writer_memory0_dat_r = mem_1[memadr_6];
assign main_sram0_dat_r0 = mem_1[memadr_7];

reg [31:0] mem_2[0:381];
reg [8:0] memadr_8;
reg [8:0] memadr_9;
always @(posedge sys_clk) begin
	if (main_writer_memory1_we)
		mem_2[main_writer_memory1_adr] <= main_writer_memory1_dat_w;
	memadr_8 <= main_writer_memory1_adr;
end

always @(posedge sys_clk) begin
	memadr_9 <= main_sram1_adr0;
end

assign main_writer_memory1_dat_r = mem_2[memadr_8];
assign main_sram1_dat_r0 = mem_2[memadr_9];

reg [31:0] mem_3[0:381];
reg [8:0] memadr_10;
reg [8:0] memadr_11;
always @(posedge sys_clk) begin
	if (main_writer_memory2_we)
		mem_3[main_writer_memory2_adr] <= main_writer_memory2_dat_w;
	memadr_10 <= main_writer_memory2_adr;
end

always @(posedge sys_clk) begin
	memadr_11 <= main_sram2_adr0;
end

assign main_writer_memory2_dat_r = mem_3[memadr_10];
assign main_sram2_dat_r0 = mem_3[memadr_11];

reg [31:0] mem_4[0:381];
reg [8:0] memadr_12;
reg [8:0] memadr_13;
always @(posedge sys_clk) begin
	if (main_writer_memory3_we)
		mem_4[main_writer_memory3_adr] <= main_writer_memory3_dat_w;
	memadr_12 <= main_writer_memory3_adr;
end

always @(posedge sys_clk) begin
	memadr_13 <= main_sram3_adr0;
end

assign main_writer_memory3_dat_r = mem_4[memadr_12];
assign main_sram3_dat_r0 = mem_4[memadr_13];

reg [13:0] storage_6[0:3];
reg [13:0] memdat_4;
always @(posedge sys_clk) begin
	if (main_reader_fifo_wrport_we)
		storage_6[main_reader_fifo_wrport_adr] <= main_reader_fifo_wrport_dat_w;
	memdat_4 <= storage_6[main_reader_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
end

assign main_reader_fifo_wrport_dat_r = memdat_4;
assign main_reader_fifo_rdport_dat_r = storage_6[main_reader_fifo_rdport_adr];

mor1kx #(
	.DBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.FEATURE_ADDC("ENABLED"),
	.FEATURE_CMOV("ENABLED"),
	.FEATURE_DATACACHE("ENABLED"),
	.FEATURE_FFL1("ENABLED"),
	.FEATURE_INSTRUCTIONCACHE("ENABLED"),
	.FEATURE_OVERFLOW("NONE"),
	.FEATURE_RANGE("NONE"),
	.FEATURE_SYSCALL("NONE"),
	.FEATURE_TIMER("NONE"),
	.FEATURE_TRAP("NONE"),
	.IBUS_WB_TYPE("B3_REGISTERED_FEEDBACK"),
	.OPTION_CPU0("CAPPUCCINO"),
	.OPTION_DCACHE_BLOCK_WIDTH(3'd4),
	.OPTION_DCACHE_LIMIT_WIDTH(5'd31),
	.OPTION_DCACHE_SET_WIDTH(4'd8),
	.OPTION_DCACHE_WAYS(1'd1),
	.OPTION_ICACHE_BLOCK_WIDTH(3'd4),
	.OPTION_ICACHE_LIMIT_WIDTH(5'd31),
	.OPTION_ICACHE_SET_WIDTH(4'd8),
	.OPTION_ICACHE_WAYS(1'd1),
	.OPTION_PIC_TRIGGER("LEVEL"),
	.OPTION_RESET_PC(31'd1082130432)
) mor1kx_1 (
	.clk(sys_kernel_clk),
	.dwbm_ack_i(main_kernel_cpu_dbus_ack),
	.dwbm_dat_i(main_kernel_cpu_dbus_dat_r),
	.dwbm_err_i(main_kernel_cpu_dbus_err),
	.dwbm_rty_i(1'd0),
	.irq_i(main_kernel_cpu_interrupt),
	.iwbm_ack_i(main_kernel_cpu_ibus_ack),
	.iwbm_dat_i(main_kernel_cpu_ibus_dat_r),
	.iwbm_err_i(main_kernel_cpu_ibus_err),
	.iwbm_rty_i(1'd0),
	.rst(sys_kernel_rst),
	.dwbm_adr_o(main_kernel_cpu_d_adr_o),
	.dwbm_bte_o(main_kernel_cpu_dbus_bte),
	.dwbm_cti_o(main_kernel_cpu_dbus_cti),
	.dwbm_cyc_o(main_kernel_cpu_dbus_cyc),
	.dwbm_dat_o(main_kernel_cpu_dbus_dat_w),
	.dwbm_sel_o(main_kernel_cpu_dbus_sel),
	.dwbm_stb_o(main_kernel_cpu_dbus_stb),
	.dwbm_we_o(main_kernel_cpu_dbus_we),
	.iwbm_adr_o(main_kernel_cpu_i_adr_o),
	.iwbm_bte_o(main_kernel_cpu_ibus_bte),
	.iwbm_cti_o(main_kernel_cpu_ibus_cti),
	.iwbm_cyc_o(main_kernel_cpu_ibus_cyc),
	.iwbm_dat_o(main_kernel_cpu_ibus_dat_w),
	.iwbm_sel_o(main_kernel_cpu_ibus_sel),
	.iwbm_stb_o(main_kernel_cpu_ibus_stb),
	.iwbm_we_o(main_kernel_cpu_ibus_we)
);

reg [7:0] mem_5[0:31];
reg [4:0] memadr_14;
always @(posedge sys_clk) begin
	memadr_14 <= main_add_identifier_adr;
end

assign main_add_identifier_dat_r = mem_5[memadr_14];

initial begin
	$readmemh("mem_5.init", mem_5);
end

assign i2c_scl = main_i2c_tstriple0_oe ? main_i2c_tstriple0_o : 1'bz;
assign main_i2c_tstriple0_i = i2c_scl;

assign i2c_sda = main_i2c_tstriple1_oe ? main_i2c_tstriple1_o : 1'bz;
assign main_i2c_tstriple1_i = i2c_sda;

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_107 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x0_o[0] ^ 1'd0)),
	.D2((main_output_8x0_o[1] ^ 1'd0)),
	.D3((main_output_8x0_o[2] ^ 1'd0)),
	.D4((main_output_8x0_o[3] ^ 1'd0)),
	.D5((main_output_8x0_o[4] ^ 1'd0)),
	.D6((main_output_8x0_o[5] ^ 1'd0)),
	.D7((main_output_8x0_o[6] ^ 1'd0)),
	.D8((main_output_8x0_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x0_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x0_pad_o),
	.TQ(main_output_8x0_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_108 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x1_o[0] ^ 1'd0)),
	.D2((main_output_8x1_o[1] ^ 1'd0)),
	.D3((main_output_8x1_o[2] ^ 1'd0)),
	.D4((main_output_8x1_o[3] ^ 1'd0)),
	.D5((main_output_8x1_o[4] ^ 1'd0)),
	.D6((main_output_8x1_o[5] ^ 1'd0)),
	.D7((main_output_8x1_o[6] ^ 1'd0)),
	.D8((main_output_8x1_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x1_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x1_pad_o),
	.TQ(main_output_8x1_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_109 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x2_o[0] ^ 1'd0)),
	.D2((main_output_8x2_o[1] ^ 1'd0)),
	.D3((main_output_8x2_o[2] ^ 1'd0)),
	.D4((main_output_8x2_o[3] ^ 1'd0)),
	.D5((main_output_8x2_o[4] ^ 1'd0)),
	.D6((main_output_8x2_o[5] ^ 1'd0)),
	.D7((main_output_8x2_o[6] ^ 1'd0)),
	.D8((main_output_8x2_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x2_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x2_pad_o),
	.TQ(main_output_8x2_t_out)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_64 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x0_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x0_serdes_i1[7]),
	.Q2(main_inout_8x0_serdes_i1[6]),
	.Q3(main_inout_8x0_serdes_i1[5]),
	.Q4(main_inout_8x0_serdes_i1[4]),
	.Q5(main_inout_8x0_serdes_i1[3]),
	.Q6(main_inout_8x0_serdes_i1[2]),
	.Q7(main_inout_8x0_serdes_i1[1]),
	.Q8(main_inout_8x0_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_110 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x0_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x0_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x0_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x0_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x0_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x0_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x0_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x0_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x0_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x0_serdes_pad_o1),
	.TQ(main_inout_8x0_serdes_t_out)
);

IOBUF IOBUF_64(
	.I(main_inout_8x0_serdes_pad_o0),
	.T(main_inout_8x0_serdes_t_out),
	.IO(ttl_3),
	.O(main_inout_8x0_serdes_pad_i0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_111 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x3_o[0] ^ 1'd0)),
	.D2((main_output_8x3_o[1] ^ 1'd0)),
	.D3((main_output_8x3_o[2] ^ 1'd0)),
	.D4((main_output_8x3_o[3] ^ 1'd0)),
	.D5((main_output_8x3_o[4] ^ 1'd0)),
	.D6((main_output_8x3_o[5] ^ 1'd0)),
	.D7((main_output_8x3_o[6] ^ 1'd0)),
	.D8((main_output_8x3_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x3_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x3_pad_o),
	.TQ(main_output_8x3_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_112 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x4_o[0] ^ 1'd0)),
	.D2((main_output_8x4_o[1] ^ 1'd0)),
	.D3((main_output_8x4_o[2] ^ 1'd0)),
	.D4((main_output_8x4_o[3] ^ 1'd0)),
	.D5((main_output_8x4_o[4] ^ 1'd0)),
	.D6((main_output_8x4_o[5] ^ 1'd0)),
	.D7((main_output_8x4_o[6] ^ 1'd0)),
	.D8((main_output_8x4_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x4_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x4_pad_o),
	.TQ(main_output_8x4_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_113 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x5_o[0] ^ 1'd0)),
	.D2((main_output_8x5_o[1] ^ 1'd0)),
	.D3((main_output_8x5_o[2] ^ 1'd0)),
	.D4((main_output_8x5_o[3] ^ 1'd0)),
	.D5((main_output_8x5_o[4] ^ 1'd0)),
	.D6((main_output_8x5_o[5] ^ 1'd0)),
	.D7((main_output_8x5_o[6] ^ 1'd0)),
	.D8((main_output_8x5_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x5_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x5_pad_o),
	.TQ(main_output_8x5_t_out)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_65 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x1_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x1_serdes_i1[7]),
	.Q2(main_inout_8x1_serdes_i1[6]),
	.Q3(main_inout_8x1_serdes_i1[5]),
	.Q4(main_inout_8x1_serdes_i1[4]),
	.Q5(main_inout_8x1_serdes_i1[3]),
	.Q6(main_inout_8x1_serdes_i1[2]),
	.Q7(main_inout_8x1_serdes_i1[1]),
	.Q8(main_inout_8x1_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_114 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x1_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x1_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x1_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x1_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x1_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x1_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x1_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x1_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x1_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x1_serdes_pad_o1),
	.TQ(main_inout_8x1_serdes_t_out)
);

IOBUF IOBUF_65(
	.I(main_inout_8x1_serdes_pad_o0),
	.T(main_inout_8x1_serdes_t_out),
	.IO(ttl_7),
	.O(main_inout_8x1_serdes_pad_i0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_115 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x6_o[0] ^ 1'd0)),
	.D2((main_output_8x6_o[1] ^ 1'd0)),
	.D3((main_output_8x6_o[2] ^ 1'd0)),
	.D4((main_output_8x6_o[3] ^ 1'd0)),
	.D5((main_output_8x6_o[4] ^ 1'd0)),
	.D6((main_output_8x6_o[5] ^ 1'd0)),
	.D7((main_output_8x6_o[6] ^ 1'd0)),
	.D8((main_output_8x6_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x6_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x6_pad_o),
	.TQ(main_output_8x6_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_116 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x7_o[0] ^ 1'd0)),
	.D2((main_output_8x7_o[1] ^ 1'd0)),
	.D3((main_output_8x7_o[2] ^ 1'd0)),
	.D4((main_output_8x7_o[3] ^ 1'd0)),
	.D5((main_output_8x7_o[4] ^ 1'd0)),
	.D6((main_output_8x7_o[5] ^ 1'd0)),
	.D7((main_output_8x7_o[6] ^ 1'd0)),
	.D8((main_output_8x7_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x7_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x7_pad_o),
	.TQ(main_output_8x7_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_117 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x8_o[0] ^ 1'd0)),
	.D2((main_output_8x8_o[1] ^ 1'd0)),
	.D3((main_output_8x8_o[2] ^ 1'd0)),
	.D4((main_output_8x8_o[3] ^ 1'd0)),
	.D5((main_output_8x8_o[4] ^ 1'd0)),
	.D6((main_output_8x8_o[5] ^ 1'd0)),
	.D7((main_output_8x8_o[6] ^ 1'd0)),
	.D8((main_output_8x8_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x8_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x8_pad_o),
	.TQ(main_output_8x8_t_out)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_66 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x2_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x2_serdes_i1[7]),
	.Q2(main_inout_8x2_serdes_i1[6]),
	.Q3(main_inout_8x2_serdes_i1[5]),
	.Q4(main_inout_8x2_serdes_i1[4]),
	.Q5(main_inout_8x2_serdes_i1[3]),
	.Q6(main_inout_8x2_serdes_i1[2]),
	.Q7(main_inout_8x2_serdes_i1[1]),
	.Q8(main_inout_8x2_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_118 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x2_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x2_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x2_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x2_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x2_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x2_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x2_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x2_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x2_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x2_serdes_pad_o1),
	.TQ(main_inout_8x2_serdes_t_out)
);

IOBUF IOBUF_66(
	.I(main_inout_8x2_serdes_pad_o0),
	.T(main_inout_8x2_serdes_t_out),
	.IO(ttl_11),
	.O(main_inout_8x2_serdes_pad_i0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_119 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x9_o[0] ^ 1'd0)),
	.D2((main_output_8x9_o[1] ^ 1'd0)),
	.D3((main_output_8x9_o[2] ^ 1'd0)),
	.D4((main_output_8x9_o[3] ^ 1'd0)),
	.D5((main_output_8x9_o[4] ^ 1'd0)),
	.D6((main_output_8x9_o[5] ^ 1'd0)),
	.D7((main_output_8x9_o[6] ^ 1'd0)),
	.D8((main_output_8x9_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x9_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x9_pad_o),
	.TQ(main_output_8x9_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_120 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x10_o[0] ^ 1'd0)),
	.D2((main_output_8x10_o[1] ^ 1'd0)),
	.D3((main_output_8x10_o[2] ^ 1'd0)),
	.D4((main_output_8x10_o[3] ^ 1'd0)),
	.D5((main_output_8x10_o[4] ^ 1'd0)),
	.D6((main_output_8x10_o[5] ^ 1'd0)),
	.D7((main_output_8x10_o[6] ^ 1'd0)),
	.D8((main_output_8x10_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x10_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x10_pad_o),
	.TQ(main_output_8x10_t_out)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_121 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_output_8x11_o[0] ^ 1'd0)),
	.D2((main_output_8x11_o[1] ^ 1'd0)),
	.D3((main_output_8x11_o[2] ^ 1'd0)),
	.D4((main_output_8x11_o[3] ^ 1'd0)),
	.D5((main_output_8x11_o[4] ^ 1'd0)),
	.D6((main_output_8x11_o[5] ^ 1'd0)),
	.D7((main_output_8x11_o[6] ^ 1'd0)),
	.D8((main_output_8x11_o[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_output_8x11_t_in),
	.TCE(1'd1),
	.OQ(main_output_8x11_pad_o),
	.TQ(main_output_8x11_t_out)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_67 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x3_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x3_serdes_i1[7]),
	.Q2(main_inout_8x3_serdes_i1[6]),
	.Q3(main_inout_8x3_serdes_i1[5]),
	.Q4(main_inout_8x3_serdes_i1[4]),
	.Q5(main_inout_8x3_serdes_i1[3]),
	.Q6(main_inout_8x3_serdes_i1[2]),
	.Q7(main_inout_8x3_serdes_i1[1]),
	.Q8(main_inout_8x3_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_122 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x3_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x3_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x3_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x3_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x3_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x3_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x3_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x3_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x3_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x3_serdes_pad_o1),
	.TQ(main_inout_8x3_serdes_t_out)
);

IOBUF IOBUF_67(
	.I(main_inout_8x3_serdes_pad_o0),
	.T(main_inout_8x3_serdes_t_out),
	.IO(ttl_15),
	.O(main_inout_8x3_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_68 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x4_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x4_serdes_i1[7]),
	.Q2(main_inout_8x4_serdes_i1[6]),
	.Q3(main_inout_8x4_serdes_i1[5]),
	.Q4(main_inout_8x4_serdes_i1[4]),
	.Q5(main_inout_8x4_serdes_i1[3]),
	.Q6(main_inout_8x4_serdes_i1[2]),
	.Q7(main_inout_8x4_serdes_i1[1]),
	.Q8(main_inout_8x4_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_123 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x4_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x4_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x4_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x4_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x4_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x4_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x4_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x4_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x4_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x4_serdes_pad_o1),
	.TQ(main_inout_8x4_serdes_t_out)
);

IOBUF IOBUF_68(
	.I(main_inout_8x4_serdes_pad_o0),
	.T(main_inout_8x4_serdes_t_out),
	.IO(pmt),
	.O(main_inout_8x4_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_69 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x5_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x5_serdes_i1[7]),
	.Q2(main_inout_8x5_serdes_i1[6]),
	.Q3(main_inout_8x5_serdes_i1[5]),
	.Q4(main_inout_8x5_serdes_i1[4]),
	.Q5(main_inout_8x5_serdes_i1[3]),
	.Q6(main_inout_8x5_serdes_i1[2]),
	.Q7(main_inout_8x5_serdes_i1[1]),
	.Q8(main_inout_8x5_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_124 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x5_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x5_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x5_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x5_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x5_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x5_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x5_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x5_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x5_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x5_serdes_pad_o1),
	.TQ(main_inout_8x5_serdes_t_out)
);

IOBUF IOBUF_69(
	.I(main_inout_8x5_serdes_pad_o0),
	.T(main_inout_8x5_serdes_t_out),
	.IO(pmt_1),
	.O(main_inout_8x5_serdes_pad_i0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.NUM_CE(1'd1)
) ISERDESE2_70 (
	.CE1(1'd1),
	.CLK(rtiox4_clk),
	.CLKB((~rtiox4_clk)),
	.CLKDIV(rio_phy_clk),
	.D(main_inout_8x6_serdes_pad_i1),
	.RST(rio_phy_rst),
	.Q1(main_inout_8x6_serdes_i1[7]),
	.Q2(main_inout_8x6_serdes_i1[6]),
	.Q3(main_inout_8x6_serdes_i1[5]),
	.Q4(main_inout_8x6_serdes_i1[4]),
	.Q5(main_inout_8x6_serdes_i1[3]),
	.Q6(main_inout_8x6_serdes_i1[2]),
	.Q7(main_inout_8x6_serdes_i1[1]),
	.Q8(main_inout_8x6_serdes_i1[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.INIT_OQ(1'd0),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_125 (
	.CLK(rtiox4_clk),
	.CLKDIV(rio_phy_clk),
	.D1((main_inout_8x6_serdes_o1[0] ^ 1'd0)),
	.D2((main_inout_8x6_serdes_o1[1] ^ 1'd0)),
	.D3((main_inout_8x6_serdes_o1[2] ^ 1'd0)),
	.D4((main_inout_8x6_serdes_o1[3] ^ 1'd0)),
	.D5((main_inout_8x6_serdes_o1[4] ^ 1'd0)),
	.D6((main_inout_8x6_serdes_o1[5] ^ 1'd0)),
	.D7((main_inout_8x6_serdes_o1[6] ^ 1'd0)),
	.D8((main_inout_8x6_serdes_o1[7] ^ 1'd0)),
	.OCE(1'd1),
	.RST(rio_phy_rst),
	.T1(main_inout_8x6_serdes_t_in),
	.TCE(1'd1),
	.OQ(main_inout_8x6_serdes_pad_o1),
	.TQ(main_inout_8x6_serdes_t_out)
);

IOBUF IOBUF_70(
	.I(main_inout_8x6_serdes_pad_o0),
	.T(main_inout_8x6_serdes_t_out),
	.IO(user_sma_gpio_n_33),
	.O(main_inout_8x6_serdes_pad_i0)
);

assign ams101_dac_cs_n = main_spimaster0_interface_cs_oe ? main_spimaster0_interface_cs_o : 1'bz;
assign main_spimaster0_interface_cs_i = ams101_dac_cs_n;

assign ams101_dac_clk = main_spimaster0_interface_clk_oe ? main_spimaster0_interface_clk_o : 1'bz;
assign main_spimaster0_interface_clk_i = ams101_dac_clk;

assign ams101_dac_mosi = main_spimaster0_interface_mosi_oe ? main_spimaster0_interface_mosi_o : 1'bz;
assign main_spimaster0_interface_mosi_i = ams101_dac_mosi;

assign spi_cs_n = main_spimaster1_interface_cs_oe ? main_spimaster1_interface_cs_o : 1'bz;
assign main_spimaster1_interface_cs_i = spi_cs_n;

assign spi_clk = main_spimaster1_interface_clk_oe ? main_spimaster1_interface_clk_o : 1'bz;
assign main_spimaster1_interface_clk_i = spi_clk;

assign spi_mosi = main_spimaster1_interface_mosi_oe ? main_spimaster1_interface_mosi_o : 1'bz;
assign main_spimaster1_interface_mosi_i = spi_mosi;

assign spi_miso = main_spimaster1_interface_miso_oe ? main_spimaster1_interface_miso_o : 1'bz;
assign main_spimaster1_interface_miso_i = spi_miso;

assign spi_cs_n_1 = main_spimaster2_interface_cs_oe ? main_spimaster2_interface_cs_o : 1'bz;
assign main_spimaster2_interface_cs_i = spi_cs_n_1;

assign spi_clk_1 = main_spimaster2_interface_clk_oe ? main_spimaster2_interface_clk_o : 1'bz;
assign main_spimaster2_interface_clk_i = spi_clk_1;

assign spi_mosi_1 = main_spimaster2_interface_mosi_oe ? main_spimaster2_interface_mosi_o : 1'bz;
assign main_spimaster2_interface_mosi_i = spi_mosi_1;

assign spi_miso_1 = main_spimaster2_interface_miso_oe ? main_spimaster2_interface_miso_o : 1'bz;
assign main_spimaster2_interface_miso_i = spi_miso_1;

assign spi_cs_n_2 = main_spimaster3_interface_cs_oe ? main_spimaster3_interface_cs_o : 1'bz;
assign main_spimaster3_interface_cs_i = spi_cs_n_2;

assign spi_clk_2 = main_spimaster3_interface_clk_oe ? main_spimaster3_interface_clk_o : 1'bz;
assign main_spimaster3_interface_clk_i = spi_clk_2;

assign spi_mosi_2 = main_spimaster3_interface_mosi_oe ? main_spimaster3_interface_mosi_o : 1'bz;
assign main_spimaster3_interface_mosi_i = spi_mosi_2;

assign spi_miso_2 = main_spimaster3_interface_miso_oe ? main_spimaster3_interface_miso_o : 1'bz;
assign main_spimaster3_interface_miso_i = spi_miso_2;

assign sdcard_spi_33_cs_n = main_spimaster4_interface_cs_oe ? main_spimaster4_interface_cs_o : 1'bz;
assign main_spimaster4_interface_cs_i = sdcard_spi_33_cs_n;

assign sdcard_spi_33_clk = main_spimaster4_interface_clk_oe ? main_spimaster4_interface_clk_o : 1'bz;
assign main_spimaster4_interface_clk_i = sdcard_spi_33_clk;

assign sdcard_spi_33_mosi = main_spimaster4_interface_mosi_oe ? main_spimaster4_interface_mosi_o : 1'bz;
assign main_spimaster4_interface_mosi_i = sdcard_spi_33_mosi;

assign sdcard_spi_33_miso = main_spimaster4_interface_miso_oe ? main_spimaster4_interface_miso_o : 1'bz;
assign main_spimaster4_interface_miso_i = sdcard_spi_33_miso;

assign dds_d = main_ad9914_oe ? main_ad9914_o : 16'bz;
assign main_ad9914_i = dds_d;

IBUFDS IBUFDS_1(
	.I(user_sma_clock_p),
	.IB(user_sma_clock_n),
	.O(main_rtio_crg_rtio_external_clk)
);

PLLE2_ADV #(
	.CLKFBOUT_MULT(4'd8),
	.CLKIN1_PERIOD(8.0),
	.CLKIN2_PERIOD(8.0),
	.CLKOUT0_DIVIDE(2'd2),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd5),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_ADV (
	.CLKFBIN(rtio_clk),
	.CLKIN1(sys_clk),
	.CLKIN2(main_rtio_crg_rtio_external_clk),
	.CLKINSEL((~main_rtio_crg_clock_sel_storage)),
	.RST(main_rtio_crg_pll_reset_storage),
	.CLKFBOUT(main_rtio_crg_rtio_clk),
	.CLKOUT0(main_rtio_crg_rtiox4_clk),
	.CLKOUT1(main_rtio_crg_ext_clkout_clk),
	.LOCKED(main_rtio_crg_pll_locked)
);

BUFG BUFG_3(
	.I(main_rtio_crg_rtio_clk),
	.O(rtio_clk)
);

BUFG BUFG_4(
	.I(main_rtio_crg_rtiox4_clk),
	.O(rtiox4_clk)
);

BUFG BUFG_5(
	.I(main_rtio_crg_ext_clkout_clk),
	.O(ext_clkout_clk)
);

reg [13:0] latency_compensation[0:28];
reg [4:0] memadr_15;
always @(posedge rsys_clk) begin
	memadr_15 <= main_rtio_core_outputs_lanedistributor_adr;
end

assign main_rtio_core_outputs_lanedistributor_dat_r = latency_compensation[memadr_15];

initial begin
	$readmemh("latency_compensation.init", latency_compensation);
end

reg [120:0] storage_7[0:127];
reg [6:0] memadr_16;
reg [6:0] memadr_17;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered0_wrport_we)
		storage_7[main_rtio_core_outputs_asyncfifobuffered0_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_w;
	memadr_16 <= main_rtio_core_outputs_asyncfifobuffered0_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_17 <= main_rtio_core_outputs_asyncfifobuffered0_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered0_wrport_dat_r = storage_7[memadr_16];
assign main_rtio_core_outputs_asyncfifobuffered0_rdport_dat_r = storage_7[memadr_17];

reg [120:0] storage_8[0:127];
reg [6:0] memadr_18;
reg [6:0] memadr_19;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered1_wrport_we)
		storage_8[main_rtio_core_outputs_asyncfifobuffered1_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_w;
	memadr_18 <= main_rtio_core_outputs_asyncfifobuffered1_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_19 <= main_rtio_core_outputs_asyncfifobuffered1_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered1_wrport_dat_r = storage_8[memadr_18];
assign main_rtio_core_outputs_asyncfifobuffered1_rdport_dat_r = storage_8[memadr_19];

reg [120:0] storage_9[0:127];
reg [6:0] memadr_20;
reg [6:0] memadr_21;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered2_wrport_we)
		storage_9[main_rtio_core_outputs_asyncfifobuffered2_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_w;
	memadr_20 <= main_rtio_core_outputs_asyncfifobuffered2_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_21 <= main_rtio_core_outputs_asyncfifobuffered2_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered2_wrport_dat_r = storage_9[memadr_20];
assign main_rtio_core_outputs_asyncfifobuffered2_rdport_dat_r = storage_9[memadr_21];

reg [120:0] storage_10[0:127];
reg [6:0] memadr_22;
reg [6:0] memadr_23;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered3_wrport_we)
		storage_10[main_rtio_core_outputs_asyncfifobuffered3_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_w;
	memadr_22 <= main_rtio_core_outputs_asyncfifobuffered3_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_23 <= main_rtio_core_outputs_asyncfifobuffered3_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered3_wrport_dat_r = storage_10[memadr_22];
assign main_rtio_core_outputs_asyncfifobuffered3_rdport_dat_r = storage_10[memadr_23];

reg [120:0] storage_11[0:127];
reg [6:0] memadr_24;
reg [6:0] memadr_25;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered4_wrport_we)
		storage_11[main_rtio_core_outputs_asyncfifobuffered4_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_w;
	memadr_24 <= main_rtio_core_outputs_asyncfifobuffered4_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_25 <= main_rtio_core_outputs_asyncfifobuffered4_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered4_wrport_dat_r = storage_11[memadr_24];
assign main_rtio_core_outputs_asyncfifobuffered4_rdport_dat_r = storage_11[memadr_25];

reg [120:0] storage_12[0:127];
reg [6:0] memadr_26;
reg [6:0] memadr_27;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered5_wrport_we)
		storage_12[main_rtio_core_outputs_asyncfifobuffered5_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_w;
	memadr_26 <= main_rtio_core_outputs_asyncfifobuffered5_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_27 <= main_rtio_core_outputs_asyncfifobuffered5_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered5_wrport_dat_r = storage_12[memadr_26];
assign main_rtio_core_outputs_asyncfifobuffered5_rdport_dat_r = storage_12[memadr_27];

reg [120:0] storage_13[0:127];
reg [6:0] memadr_28;
reg [6:0] memadr_29;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered6_wrport_we)
		storage_13[main_rtio_core_outputs_asyncfifobuffered6_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_w;
	memadr_28 <= main_rtio_core_outputs_asyncfifobuffered6_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_29 <= main_rtio_core_outputs_asyncfifobuffered6_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered6_wrport_dat_r = storage_13[memadr_28];
assign main_rtio_core_outputs_asyncfifobuffered6_rdport_dat_r = storage_13[memadr_29];

reg [120:0] storage_14[0:127];
reg [6:0] memadr_30;
reg [6:0] memadr_31;
always @(posedge rsys_clk) begin
	if (main_rtio_core_outputs_asyncfifobuffered7_wrport_we)
		storage_14[main_rtio_core_outputs_asyncfifobuffered7_wrport_adr] <= main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_w;
	memadr_30 <= main_rtio_core_outputs_asyncfifobuffered7_wrport_adr;
end

always @(posedge rio_clk) begin
	memadr_31 <= main_rtio_core_outputs_asyncfifobuffered7_rdport_adr;
end

assign main_rtio_core_outputs_asyncfifobuffered7_wrport_dat_r = storage_14[memadr_30];
assign main_rtio_core_outputs_asyncfifobuffered7_rdport_dat_r = storage_14[memadr_31];

reg [0:0] en_replaces_rom[0:28];
reg [4:0] memadr_32;
always @(posedge rio_clk) begin
	memadr_32 <= main_rtio_core_outputs_memory0_adr;
end

assign main_rtio_core_outputs_memory0_dat_r = en_replaces_rom[memadr_32];

initial begin
	$readmemh("en_replaces_rom.init", en_replaces_rom);
end

reg [0:0] en_replaces_rom_1[0:28];
reg [4:0] memadr_33;
always @(posedge rio_clk) begin
	memadr_33 <= main_rtio_core_outputs_memory1_adr;
end

assign main_rtio_core_outputs_memory1_dat_r = en_replaces_rom_1[memadr_33];

initial begin
	$readmemh("en_replaces_rom_1.init", en_replaces_rom_1);
end

reg [0:0] en_replaces_rom_2[0:28];
reg [4:0] memadr_34;
always @(posedge rio_clk) begin
	memadr_34 <= main_rtio_core_outputs_memory2_adr;
end

assign main_rtio_core_outputs_memory2_dat_r = en_replaces_rom_2[memadr_34];

initial begin
	$readmemh("en_replaces_rom_2.init", en_replaces_rom_2);
end

reg [0:0] en_replaces_rom_3[0:28];
reg [4:0] memadr_35;
always @(posedge rio_clk) begin
	memadr_35 <= main_rtio_core_outputs_memory3_adr;
end

assign main_rtio_core_outputs_memory3_dat_r = en_replaces_rom_3[memadr_35];

initial begin
	$readmemh("en_replaces_rom_3.init", en_replaces_rom_3);
end

reg [0:0] en_replaces_rom_4[0:28];
reg [4:0] memadr_36;
always @(posedge rio_clk) begin
	memadr_36 <= main_rtio_core_outputs_memory4_adr;
end

assign main_rtio_core_outputs_memory4_dat_r = en_replaces_rom_4[memadr_36];

initial begin
	$readmemh("en_replaces_rom_4.init", en_replaces_rom_4);
end

reg [0:0] en_replaces_rom_5[0:28];
reg [4:0] memadr_37;
always @(posedge rio_clk) begin
	memadr_37 <= main_rtio_core_outputs_memory5_adr;
end

assign main_rtio_core_outputs_memory5_dat_r = en_replaces_rom_5[memadr_37];

initial begin
	$readmemh("en_replaces_rom_5.init", en_replaces_rom_5);
end

reg [0:0] en_replaces_rom_6[0:28];
reg [4:0] memadr_38;
always @(posedge rio_clk) begin
	memadr_38 <= main_rtio_core_outputs_memory6_adr;
end

assign main_rtio_core_outputs_memory6_dat_r = en_replaces_rom_6[memadr_38];

initial begin
	$readmemh("en_replaces_rom_6.init", en_replaces_rom_6);
end

reg [0:0] en_replaces_rom_7[0:28];
reg [4:0] memadr_39;
always @(posedge rio_clk) begin
	memadr_39 <= main_rtio_core_outputs_memory7_adr;
end

assign main_rtio_core_outputs_memory7_dat_r = en_replaces_rom_7[memadr_39];

initial begin
	$readmemh("en_replaces_rom_7.init", en_replaces_rom_7);
end

reg [64:0] storage_15[0:511];
reg [8:0] memadr_40;
reg [8:0] memadr_41;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo0_wrport_we)
		storage_15[main_rtio_core_inputs_asyncfifo0_wrport_adr] <= main_rtio_core_inputs_asyncfifo0_wrport_dat_w;
	memadr_40 <= main_rtio_core_inputs_asyncfifo0_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_41 <= main_rtio_core_inputs_asyncfifo0_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo0_wrport_dat_r = storage_15[memadr_40];
assign main_rtio_core_inputs_asyncfifo0_rdport_dat_r = storage_15[memadr_41];

reg [64:0] storage_16[0:511];
reg [8:0] memadr_42;
reg [8:0] memadr_43;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo1_wrport_we)
		storage_16[main_rtio_core_inputs_asyncfifo1_wrport_adr] <= main_rtio_core_inputs_asyncfifo1_wrport_dat_w;
	memadr_42 <= main_rtio_core_inputs_asyncfifo1_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_43 <= main_rtio_core_inputs_asyncfifo1_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo1_wrport_dat_r = storage_16[memadr_42];
assign main_rtio_core_inputs_asyncfifo1_rdport_dat_r = storage_16[memadr_43];

reg [64:0] storage_17[0:511];
reg [8:0] memadr_44;
reg [8:0] memadr_45;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo2_wrport_we)
		storage_17[main_rtio_core_inputs_asyncfifo2_wrport_adr] <= main_rtio_core_inputs_asyncfifo2_wrport_dat_w;
	memadr_44 <= main_rtio_core_inputs_asyncfifo2_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_45 <= main_rtio_core_inputs_asyncfifo2_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo2_wrport_dat_r = storage_17[memadr_44];
assign main_rtio_core_inputs_asyncfifo2_rdport_dat_r = storage_17[memadr_45];

reg [64:0] storage_18[0:511];
reg [8:0] memadr_46;
reg [8:0] memadr_47;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo3_wrport_we)
		storage_18[main_rtio_core_inputs_asyncfifo3_wrport_adr] <= main_rtio_core_inputs_asyncfifo3_wrport_dat_w;
	memadr_46 <= main_rtio_core_inputs_asyncfifo3_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_47 <= main_rtio_core_inputs_asyncfifo3_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo3_wrport_dat_r = storage_18[memadr_46];
assign main_rtio_core_inputs_asyncfifo3_rdport_dat_r = storage_18[memadr_47];

reg [64:0] storage_19[0:511];
reg [8:0] memadr_48;
reg [8:0] memadr_49;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo4_wrport_we)
		storage_19[main_rtio_core_inputs_asyncfifo4_wrport_adr] <= main_rtio_core_inputs_asyncfifo4_wrport_dat_w;
	memadr_48 <= main_rtio_core_inputs_asyncfifo4_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_49 <= main_rtio_core_inputs_asyncfifo4_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo4_wrport_dat_r = storage_19[memadr_48];
assign main_rtio_core_inputs_asyncfifo4_rdport_dat_r = storage_19[memadr_49];

reg [64:0] storage_20[0:511];
reg [8:0] memadr_50;
reg [8:0] memadr_51;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo5_wrport_we)
		storage_20[main_rtio_core_inputs_asyncfifo5_wrport_adr] <= main_rtio_core_inputs_asyncfifo5_wrport_dat_w;
	memadr_50 <= main_rtio_core_inputs_asyncfifo5_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_51 <= main_rtio_core_inputs_asyncfifo5_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo5_wrport_dat_r = storage_20[memadr_50];
assign main_rtio_core_inputs_asyncfifo5_rdport_dat_r = storage_20[memadr_51];

reg [64:0] storage_21[0:511];
reg [8:0] memadr_52;
reg [8:0] memadr_53;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo6_wrport_we)
		storage_21[main_rtio_core_inputs_asyncfifo6_wrport_adr] <= main_rtio_core_inputs_asyncfifo6_wrport_dat_w;
	memadr_52 <= main_rtio_core_inputs_asyncfifo6_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_53 <= main_rtio_core_inputs_asyncfifo6_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo6_wrport_dat_r = storage_21[memadr_52];
assign main_rtio_core_inputs_asyncfifo6_rdport_dat_r = storage_21[memadr_53];

reg [31:0] storage_22[0:3];
reg [1:0] memadr_54;
reg [1:0] memadr_55;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo7_wrport_we)
		storage_22[main_rtio_core_inputs_asyncfifo7_wrport_adr] <= main_rtio_core_inputs_asyncfifo7_wrport_dat_w;
	memadr_54 <= main_rtio_core_inputs_asyncfifo7_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_55 <= main_rtio_core_inputs_asyncfifo7_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo7_wrport_dat_r = storage_22[memadr_54];
assign main_rtio_core_inputs_asyncfifo7_rdport_dat_r = storage_22[memadr_55];

reg [31:0] storage_23[0:127];
reg [6:0] memadr_56;
reg [6:0] memadr_57;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo8_wrport_we)
		storage_23[main_rtio_core_inputs_asyncfifo8_wrport_adr] <= main_rtio_core_inputs_asyncfifo8_wrport_dat_w;
	memadr_56 <= main_rtio_core_inputs_asyncfifo8_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_57 <= main_rtio_core_inputs_asyncfifo8_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo8_wrport_dat_r = storage_23[memadr_56];
assign main_rtio_core_inputs_asyncfifo8_rdport_dat_r = storage_23[memadr_57];

reg [31:0] storage_24[0:127];
reg [6:0] memadr_58;
reg [6:0] memadr_59;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo9_wrport_we)
		storage_24[main_rtio_core_inputs_asyncfifo9_wrport_adr] <= main_rtio_core_inputs_asyncfifo9_wrport_dat_w;
	memadr_58 <= main_rtio_core_inputs_asyncfifo9_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_59 <= main_rtio_core_inputs_asyncfifo9_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo9_wrport_dat_r = storage_24[memadr_58];
assign main_rtio_core_inputs_asyncfifo9_rdport_dat_r = storage_24[memadr_59];

reg [31:0] storage_25[0:127];
reg [6:0] memadr_60;
reg [6:0] memadr_61;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo10_wrport_we)
		storage_25[main_rtio_core_inputs_asyncfifo10_wrport_adr] <= main_rtio_core_inputs_asyncfifo10_wrport_dat_w;
	memadr_60 <= main_rtio_core_inputs_asyncfifo10_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_61 <= main_rtio_core_inputs_asyncfifo10_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo10_wrport_dat_r = storage_25[memadr_60];
assign main_rtio_core_inputs_asyncfifo10_rdport_dat_r = storage_25[memadr_61];

reg [31:0] storage_26[0:3];
reg [1:0] memadr_62;
reg [1:0] memadr_63;
always @(posedge rio_clk) begin
	if (main_rtio_core_inputs_asyncfifo11_wrport_we)
		storage_26[main_rtio_core_inputs_asyncfifo11_wrport_adr] <= main_rtio_core_inputs_asyncfifo11_wrport_dat_w;
	memadr_62 <= main_rtio_core_inputs_asyncfifo11_wrport_adr;
end

always @(posedge rsys_clk) begin
	memadr_63 <= main_rtio_core_inputs_asyncfifo11_rdport_adr;
end

assign main_rtio_core_inputs_asyncfifo11_wrport_dat_r = storage_26[memadr_62];
assign main_rtio_core_inputs_asyncfifo11_rdport_dat_r = storage_26[memadr_63];

reg [256:0] storage_27[0:127];
reg [256:0] memdat_5;
reg [256:0] memdat_6;
always @(posedge sys_clk) begin
	if (main_rtio_analyzer_fifo_wrport_we)
		storage_27[main_rtio_analyzer_fifo_wrport_adr] <= main_rtio_analyzer_fifo_wrport_dat_w;
	memdat_5 <= storage_27[main_rtio_analyzer_fifo_wrport_adr];
end

always @(posedge sys_clk) begin
	if (main_rtio_analyzer_fifo_rdport_re)
		memdat_6 <= storage_27[main_rtio_analyzer_fifo_rdport_adr];
end

assign main_rtio_analyzer_fifo_wrport_dat_r = memdat_5;
assign main_rtio_analyzer_fifo_rdport_dat_r = memdat_6;

reg [7:0] data_mem_grain0[0:2047];
reg [10:0] memadr_64;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[0])
		data_mem_grain0[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[7:0];
	memadr_64 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[7:0] = data_mem_grain0[memadr_64];

reg [7:0] data_mem_grain1[0:2047];
reg [10:0] memadr_65;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[1])
		data_mem_grain1[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[15:8];
	memadr_65 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[15:8] = data_mem_grain1[memadr_65];

reg [7:0] data_mem_grain2[0:2047];
reg [10:0] memadr_66;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[2])
		data_mem_grain2[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[23:16];
	memadr_66 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[23:16] = data_mem_grain2[memadr_66];

reg [7:0] data_mem_grain3[0:2047];
reg [10:0] memadr_67;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[3])
		data_mem_grain3[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[31:24];
	memadr_67 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[31:24] = data_mem_grain3[memadr_67];

reg [7:0] data_mem_grain4[0:2047];
reg [10:0] memadr_68;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[4])
		data_mem_grain4[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[39:32];
	memadr_68 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[39:32] = data_mem_grain4[memadr_68];

reg [7:0] data_mem_grain5[0:2047];
reg [10:0] memadr_69;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[5])
		data_mem_grain5[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[47:40];
	memadr_69 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[47:40] = data_mem_grain5[memadr_69];

reg [7:0] data_mem_grain6[0:2047];
reg [10:0] memadr_70;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[6])
		data_mem_grain6[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[55:48];
	memadr_70 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[55:48] = data_mem_grain6[memadr_70];

reg [7:0] data_mem_grain7[0:2047];
reg [10:0] memadr_71;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[7])
		data_mem_grain7[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[63:56];
	memadr_71 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[63:56] = data_mem_grain7[memadr_71];

reg [7:0] data_mem_grain8[0:2047];
reg [10:0] memadr_72;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[8])
		data_mem_grain8[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[71:64];
	memadr_72 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[71:64] = data_mem_grain8[memadr_72];

reg [7:0] data_mem_grain9[0:2047];
reg [10:0] memadr_73;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[9])
		data_mem_grain9[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[79:72];
	memadr_73 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[79:72] = data_mem_grain9[memadr_73];

reg [7:0] data_mem_grain10[0:2047];
reg [10:0] memadr_74;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[10])
		data_mem_grain10[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[87:80];
	memadr_74 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[87:80] = data_mem_grain10[memadr_74];

reg [7:0] data_mem_grain11[0:2047];
reg [10:0] memadr_75;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[11])
		data_mem_grain11[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[95:88];
	memadr_75 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[95:88] = data_mem_grain11[memadr_75];

reg [7:0] data_mem_grain12[0:2047];
reg [10:0] memadr_76;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[12])
		data_mem_grain12[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[103:96];
	memadr_76 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[103:96] = data_mem_grain12[memadr_76];

reg [7:0] data_mem_grain13[0:2047];
reg [10:0] memadr_77;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[13])
		data_mem_grain13[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[111:104];
	memadr_77 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[111:104] = data_mem_grain13[memadr_77];

reg [7:0] data_mem_grain14[0:2047];
reg [10:0] memadr_78;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[14])
		data_mem_grain14[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[119:112];
	memadr_78 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[119:112] = data_mem_grain14[memadr_78];

reg [7:0] data_mem_grain15[0:2047];
reg [10:0] memadr_79;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[15])
		data_mem_grain15[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[127:120];
	memadr_79 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[127:120] = data_mem_grain15[memadr_79];

reg [7:0] data_mem_grain16[0:2047];
reg [10:0] memadr_80;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[16])
		data_mem_grain16[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[135:128];
	memadr_80 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[135:128] = data_mem_grain16[memadr_80];

reg [7:0] data_mem_grain17[0:2047];
reg [10:0] memadr_81;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[17])
		data_mem_grain17[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[143:136];
	memadr_81 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[143:136] = data_mem_grain17[memadr_81];

reg [7:0] data_mem_grain18[0:2047];
reg [10:0] memadr_82;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[18])
		data_mem_grain18[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[151:144];
	memadr_82 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[151:144] = data_mem_grain18[memadr_82];

reg [7:0] data_mem_grain19[0:2047];
reg [10:0] memadr_83;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[19])
		data_mem_grain19[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[159:152];
	memadr_83 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[159:152] = data_mem_grain19[memadr_83];

reg [7:0] data_mem_grain20[0:2047];
reg [10:0] memadr_84;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[20])
		data_mem_grain20[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[167:160];
	memadr_84 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[167:160] = data_mem_grain20[memadr_84];

reg [7:0] data_mem_grain21[0:2047];
reg [10:0] memadr_85;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[21])
		data_mem_grain21[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[175:168];
	memadr_85 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[175:168] = data_mem_grain21[memadr_85];

reg [7:0] data_mem_grain22[0:2047];
reg [10:0] memadr_86;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[22])
		data_mem_grain22[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[183:176];
	memadr_86 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[183:176] = data_mem_grain22[memadr_86];

reg [7:0] data_mem_grain23[0:2047];
reg [10:0] memadr_87;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[23])
		data_mem_grain23[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[191:184];
	memadr_87 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[191:184] = data_mem_grain23[memadr_87];

reg [7:0] data_mem_grain24[0:2047];
reg [10:0] memadr_88;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[24])
		data_mem_grain24[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[199:192];
	memadr_88 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[199:192] = data_mem_grain24[memadr_88];

reg [7:0] data_mem_grain25[0:2047];
reg [10:0] memadr_89;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[25])
		data_mem_grain25[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[207:200];
	memadr_89 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[207:200] = data_mem_grain25[memadr_89];

reg [7:0] data_mem_grain26[0:2047];
reg [10:0] memadr_90;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[26])
		data_mem_grain26[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[215:208];
	memadr_90 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[215:208] = data_mem_grain26[memadr_90];

reg [7:0] data_mem_grain27[0:2047];
reg [10:0] memadr_91;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[27])
		data_mem_grain27[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[223:216];
	memadr_91 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[223:216] = data_mem_grain27[memadr_91];

reg [7:0] data_mem_grain28[0:2047];
reg [10:0] memadr_92;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[28])
		data_mem_grain28[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[231:224];
	memadr_92 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[231:224] = data_mem_grain28[memadr_92];

reg [7:0] data_mem_grain29[0:2047];
reg [10:0] memadr_93;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[29])
		data_mem_grain29[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[239:232];
	memadr_93 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[239:232] = data_mem_grain29[memadr_93];

reg [7:0] data_mem_grain30[0:2047];
reg [10:0] memadr_94;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[30])
		data_mem_grain30[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[247:240];
	memadr_94 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[247:240] = data_mem_grain30[memadr_94];

reg [7:0] data_mem_grain31[0:2047];
reg [10:0] memadr_95;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[31])
		data_mem_grain31[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[255:248];
	memadr_95 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[255:248] = data_mem_grain31[memadr_95];

reg [7:0] data_mem_grain32[0:2047];
reg [10:0] memadr_96;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[32])
		data_mem_grain32[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[263:256];
	memadr_96 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[263:256] = data_mem_grain32[memadr_96];

reg [7:0] data_mem_grain33[0:2047];
reg [10:0] memadr_97;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[33])
		data_mem_grain33[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[271:264];
	memadr_97 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[271:264] = data_mem_grain33[memadr_97];

reg [7:0] data_mem_grain34[0:2047];
reg [10:0] memadr_98;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[34])
		data_mem_grain34[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[279:272];
	memadr_98 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[279:272] = data_mem_grain34[memadr_98];

reg [7:0] data_mem_grain35[0:2047];
reg [10:0] memadr_99;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[35])
		data_mem_grain35[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[287:280];
	memadr_99 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[287:280] = data_mem_grain35[memadr_99];

reg [7:0] data_mem_grain36[0:2047];
reg [10:0] memadr_100;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[36])
		data_mem_grain36[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[295:288];
	memadr_100 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[295:288] = data_mem_grain36[memadr_100];

reg [7:0] data_mem_grain37[0:2047];
reg [10:0] memadr_101;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[37])
		data_mem_grain37[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[303:296];
	memadr_101 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[303:296] = data_mem_grain37[memadr_101];

reg [7:0] data_mem_grain38[0:2047];
reg [10:0] memadr_102;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[38])
		data_mem_grain38[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[311:304];
	memadr_102 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[311:304] = data_mem_grain38[memadr_102];

reg [7:0] data_mem_grain39[0:2047];
reg [10:0] memadr_103;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[39])
		data_mem_grain39[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[319:312];
	memadr_103 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[319:312] = data_mem_grain39[memadr_103];

reg [7:0] data_mem_grain40[0:2047];
reg [10:0] memadr_104;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[40])
		data_mem_grain40[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[327:320];
	memadr_104 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[327:320] = data_mem_grain40[memadr_104];

reg [7:0] data_mem_grain41[0:2047];
reg [10:0] memadr_105;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[41])
		data_mem_grain41[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[335:328];
	memadr_105 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[335:328] = data_mem_grain41[memadr_105];

reg [7:0] data_mem_grain42[0:2047];
reg [10:0] memadr_106;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[42])
		data_mem_grain42[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[343:336];
	memadr_106 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[343:336] = data_mem_grain42[memadr_106];

reg [7:0] data_mem_grain43[0:2047];
reg [10:0] memadr_107;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[43])
		data_mem_grain43[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[351:344];
	memadr_107 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[351:344] = data_mem_grain43[memadr_107];

reg [7:0] data_mem_grain44[0:2047];
reg [10:0] memadr_108;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[44])
		data_mem_grain44[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[359:352];
	memadr_108 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[359:352] = data_mem_grain44[memadr_108];

reg [7:0] data_mem_grain45[0:2047];
reg [10:0] memadr_109;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[45])
		data_mem_grain45[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[367:360];
	memadr_109 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[367:360] = data_mem_grain45[memadr_109];

reg [7:0] data_mem_grain46[0:2047];
reg [10:0] memadr_110;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[46])
		data_mem_grain46[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[375:368];
	memadr_110 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[375:368] = data_mem_grain46[memadr_110];

reg [7:0] data_mem_grain47[0:2047];
reg [10:0] memadr_111;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[47])
		data_mem_grain47[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[383:376];
	memadr_111 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[383:376] = data_mem_grain47[memadr_111];

reg [7:0] data_mem_grain48[0:2047];
reg [10:0] memadr_112;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[48])
		data_mem_grain48[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[391:384];
	memadr_112 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[391:384] = data_mem_grain48[memadr_112];

reg [7:0] data_mem_grain49[0:2047];
reg [10:0] memadr_113;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[49])
		data_mem_grain49[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[399:392];
	memadr_113 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[399:392] = data_mem_grain49[memadr_113];

reg [7:0] data_mem_grain50[0:2047];
reg [10:0] memadr_114;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[50])
		data_mem_grain50[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[407:400];
	memadr_114 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[407:400] = data_mem_grain50[memadr_114];

reg [7:0] data_mem_grain51[0:2047];
reg [10:0] memadr_115;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[51])
		data_mem_grain51[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[415:408];
	memadr_115 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[415:408] = data_mem_grain51[memadr_115];

reg [7:0] data_mem_grain52[0:2047];
reg [10:0] memadr_116;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[52])
		data_mem_grain52[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[423:416];
	memadr_116 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[423:416] = data_mem_grain52[memadr_116];

reg [7:0] data_mem_grain53[0:2047];
reg [10:0] memadr_117;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[53])
		data_mem_grain53[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[431:424];
	memadr_117 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[431:424] = data_mem_grain53[memadr_117];

reg [7:0] data_mem_grain54[0:2047];
reg [10:0] memadr_118;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[54])
		data_mem_grain54[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[439:432];
	memadr_118 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[439:432] = data_mem_grain54[memadr_118];

reg [7:0] data_mem_grain55[0:2047];
reg [10:0] memadr_119;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[55])
		data_mem_grain55[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[447:440];
	memadr_119 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[447:440] = data_mem_grain55[memadr_119];

reg [7:0] data_mem_grain56[0:2047];
reg [10:0] memadr_120;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[56])
		data_mem_grain56[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[455:448];
	memadr_120 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[455:448] = data_mem_grain56[memadr_120];

reg [7:0] data_mem_grain57[0:2047];
reg [10:0] memadr_121;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[57])
		data_mem_grain57[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[463:456];
	memadr_121 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[463:456] = data_mem_grain57[memadr_121];

reg [7:0] data_mem_grain58[0:2047];
reg [10:0] memadr_122;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[58])
		data_mem_grain58[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[471:464];
	memadr_122 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[471:464] = data_mem_grain58[memadr_122];

reg [7:0] data_mem_grain59[0:2047];
reg [10:0] memadr_123;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[59])
		data_mem_grain59[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[479:472];
	memadr_123 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[479:472] = data_mem_grain59[memadr_123];

reg [7:0] data_mem_grain60[0:2047];
reg [10:0] memadr_124;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[60])
		data_mem_grain60[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[487:480];
	memadr_124 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[487:480] = data_mem_grain60[memadr_124];

reg [7:0] data_mem_grain61[0:2047];
reg [10:0] memadr_125;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[61])
		data_mem_grain61[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[495:488];
	memadr_125 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[495:488] = data_mem_grain61[memadr_125];

reg [7:0] data_mem_grain62[0:2047];
reg [10:0] memadr_126;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[62])
		data_mem_grain62[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[503:496];
	memadr_126 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[503:496] = data_mem_grain62[memadr_126];

reg [7:0] data_mem_grain63[0:2047];
reg [10:0] memadr_127;
always @(posedge sys_clk) begin
	if (main_nist_clock_nist_clock_data_port_we[63])
		data_mem_grain63[main_nist_clock_nist_clock_data_port_adr] <= main_nist_clock_nist_clock_data_port_dat_w[511:504];
	memadr_127 <= main_nist_clock_nist_clock_data_port_adr;
end

assign main_nist_clock_nist_clock_data_port_dat_r[511:504] = data_mem_grain63[memadr_127];

reg [7:0] mem_grain0[0:381];
reg [8:0] memadr_128;
reg [8:0] memadr_129;
always @(posedge sys_clk) begin
	memadr_128 <= main_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_sram0_we[0])
		mem_grain0[main_sram0_adr1] <= main_sram0_dat_w[7:0];
	memadr_129 <= main_sram0_adr1;
end

assign main_reader_memory0_dat_r[7:0] = mem_grain0[memadr_128];
assign main_sram0_dat_r1[7:0] = mem_grain0[memadr_129];

reg [7:0] mem_grain1[0:381];
reg [8:0] memadr_130;
reg [8:0] memadr_131;
always @(posedge sys_clk) begin
	memadr_130 <= main_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_sram0_we[1])
		mem_grain1[main_sram0_adr1] <= main_sram0_dat_w[15:8];
	memadr_131 <= main_sram0_adr1;
end

assign main_reader_memory0_dat_r[15:8] = mem_grain1[memadr_130];
assign main_sram0_dat_r1[15:8] = mem_grain1[memadr_131];

reg [7:0] mem_grain2[0:381];
reg [8:0] memadr_132;
reg [8:0] memadr_133;
always @(posedge sys_clk) begin
	memadr_132 <= main_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_sram0_we[2])
		mem_grain2[main_sram0_adr1] <= main_sram0_dat_w[23:16];
	memadr_133 <= main_sram0_adr1;
end

assign main_reader_memory0_dat_r[23:16] = mem_grain2[memadr_132];
assign main_sram0_dat_r1[23:16] = mem_grain2[memadr_133];

reg [7:0] mem_grain3[0:381];
reg [8:0] memadr_134;
reg [8:0] memadr_135;
always @(posedge sys_clk) begin
	memadr_134 <= main_reader_memory0_adr;
end

always @(posedge sys_clk) begin
	if (main_sram0_we[3])
		mem_grain3[main_sram0_adr1] <= main_sram0_dat_w[31:24];
	memadr_135 <= main_sram0_adr1;
end

assign main_reader_memory0_dat_r[31:24] = mem_grain3[memadr_134];
assign main_sram0_dat_r1[31:24] = mem_grain3[memadr_135];

reg [7:0] mem_grain0_1[0:381];
reg [8:0] memadr_136;
reg [8:0] memadr_137;
always @(posedge sys_clk) begin
	memadr_136 <= main_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_sram1_we[0])
		mem_grain0_1[main_sram1_adr1] <= main_sram1_dat_w[7:0];
	memadr_137 <= main_sram1_adr1;
end

assign main_reader_memory1_dat_r[7:0] = mem_grain0_1[memadr_136];
assign main_sram1_dat_r1[7:0] = mem_grain0_1[memadr_137];

reg [7:0] mem_grain1_1[0:381];
reg [8:0] memadr_138;
reg [8:0] memadr_139;
always @(posedge sys_clk) begin
	memadr_138 <= main_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_sram1_we[1])
		mem_grain1_1[main_sram1_adr1] <= main_sram1_dat_w[15:8];
	memadr_139 <= main_sram1_adr1;
end

assign main_reader_memory1_dat_r[15:8] = mem_grain1_1[memadr_138];
assign main_sram1_dat_r1[15:8] = mem_grain1_1[memadr_139];

reg [7:0] mem_grain2_1[0:381];
reg [8:0] memadr_140;
reg [8:0] memadr_141;
always @(posedge sys_clk) begin
	memadr_140 <= main_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_sram1_we[2])
		mem_grain2_1[main_sram1_adr1] <= main_sram1_dat_w[23:16];
	memadr_141 <= main_sram1_adr1;
end

assign main_reader_memory1_dat_r[23:16] = mem_grain2_1[memadr_140];
assign main_sram1_dat_r1[23:16] = mem_grain2_1[memadr_141];

reg [7:0] mem_grain3_1[0:381];
reg [8:0] memadr_142;
reg [8:0] memadr_143;
always @(posedge sys_clk) begin
	memadr_142 <= main_reader_memory1_adr;
end

always @(posedge sys_clk) begin
	if (main_sram1_we[3])
		mem_grain3_1[main_sram1_adr1] <= main_sram1_dat_w[31:24];
	memadr_143 <= main_sram1_adr1;
end

assign main_reader_memory1_dat_r[31:24] = mem_grain3_1[memadr_142];
assign main_sram1_dat_r1[31:24] = mem_grain3_1[memadr_143];

reg [7:0] mem_grain0_2[0:381];
reg [8:0] memadr_144;
reg [8:0] memadr_145;
always @(posedge sys_clk) begin
	memadr_144 <= main_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_sram2_we[0])
		mem_grain0_2[main_sram2_adr1] <= main_sram2_dat_w[7:0];
	memadr_145 <= main_sram2_adr1;
end

assign main_reader_memory2_dat_r[7:0] = mem_grain0_2[memadr_144];
assign main_sram2_dat_r1[7:0] = mem_grain0_2[memadr_145];

reg [7:0] mem_grain1_2[0:381];
reg [8:0] memadr_146;
reg [8:0] memadr_147;
always @(posedge sys_clk) begin
	memadr_146 <= main_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_sram2_we[1])
		mem_grain1_2[main_sram2_adr1] <= main_sram2_dat_w[15:8];
	memadr_147 <= main_sram2_adr1;
end

assign main_reader_memory2_dat_r[15:8] = mem_grain1_2[memadr_146];
assign main_sram2_dat_r1[15:8] = mem_grain1_2[memadr_147];

reg [7:0] mem_grain2_2[0:381];
reg [8:0] memadr_148;
reg [8:0] memadr_149;
always @(posedge sys_clk) begin
	memadr_148 <= main_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_sram2_we[2])
		mem_grain2_2[main_sram2_adr1] <= main_sram2_dat_w[23:16];
	memadr_149 <= main_sram2_adr1;
end

assign main_reader_memory2_dat_r[23:16] = mem_grain2_2[memadr_148];
assign main_sram2_dat_r1[23:16] = mem_grain2_2[memadr_149];

reg [7:0] mem_grain3_2[0:381];
reg [8:0] memadr_150;
reg [8:0] memadr_151;
always @(posedge sys_clk) begin
	memadr_150 <= main_reader_memory2_adr;
end

always @(posedge sys_clk) begin
	if (main_sram2_we[3])
		mem_grain3_2[main_sram2_adr1] <= main_sram2_dat_w[31:24];
	memadr_151 <= main_sram2_adr1;
end

assign main_reader_memory2_dat_r[31:24] = mem_grain3_2[memadr_150];
assign main_sram2_dat_r1[31:24] = mem_grain3_2[memadr_151];

reg [7:0] mem_grain0_3[0:381];
reg [8:0] memadr_152;
reg [8:0] memadr_153;
always @(posedge sys_clk) begin
	memadr_152 <= main_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_sram3_we[0])
		mem_grain0_3[main_sram3_adr1] <= main_sram3_dat_w[7:0];
	memadr_153 <= main_sram3_adr1;
end

assign main_reader_memory3_dat_r[7:0] = mem_grain0_3[memadr_152];
assign main_sram3_dat_r1[7:0] = mem_grain0_3[memadr_153];

reg [7:0] mem_grain1_3[0:381];
reg [8:0] memadr_154;
reg [8:0] memadr_155;
always @(posedge sys_clk) begin
	memadr_154 <= main_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_sram3_we[1])
		mem_grain1_3[main_sram3_adr1] <= main_sram3_dat_w[15:8];
	memadr_155 <= main_sram3_adr1;
end

assign main_reader_memory3_dat_r[15:8] = mem_grain1_3[memadr_154];
assign main_sram3_dat_r1[15:8] = mem_grain1_3[memadr_155];

reg [7:0] mem_grain2_3[0:381];
reg [8:0] memadr_156;
reg [8:0] memadr_157;
always @(posedge sys_clk) begin
	memadr_156 <= main_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_sram3_we[2])
		mem_grain2_3[main_sram3_adr1] <= main_sram3_dat_w[23:16];
	memadr_157 <= main_sram3_adr1;
end

assign main_reader_memory3_dat_r[23:16] = mem_grain2_3[memadr_156];
assign main_sram3_dat_r1[23:16] = mem_grain2_3[memadr_157];

reg [7:0] mem_grain3_3[0:381];
reg [8:0] memadr_158;
reg [8:0] memadr_159;
always @(posedge sys_clk) begin
	memadr_158 <= main_reader_memory3_adr;
end

always @(posedge sys_clk) begin
	if (main_sram3_we[3])
		mem_grain3_3[main_sram3_adr1] <= main_sram3_dat_w[31:24];
	memadr_159 <= main_sram3_adr1;
end

assign main_reader_memory3_dat_r[31:24] = mem_grain3_3[memadr_158];
assign main_sram3_dat_r1[31:24] = mem_grain3_3[memadr_159];

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(builder_xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(sys_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(builder_xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(clk200_rst)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(1'd1),
	.D2((main_ethphy_mode0 == 1'd1)),
	.R(1'd0),
	.S(1'd0),
	.Q(eth_clocks_gtx)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_ethphy_storage),
	.Q(builder_xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(main_ethphy_storage),
	.Q(eth_tx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_ethphy_storage),
	.Q(builder_xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(main_ethphy_storage),
	.Q(eth_rx_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl4),
	.Q(builder_xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(rtio_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl4),
	.Q(rtio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(rio_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_rtio_core_cmd_reset),
	.Q(builder_xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(rio_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(main_rtio_core_cmd_reset),
	.Q(rio_rst)
);

(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(main_rtio_core_cmd_reset_phy),
	.Q(builder_xilinxasyncresetsynchronizerimpl6_rst_meta)
);

(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(rio_phy_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl6_rst_meta),
	.PRE(main_rtio_core_cmd_reset_phy),
	.Q(rio_phy_rst)
);

endmodule
